##
## LEF for PtnCells ;
## created by Innovus v19.17-s077_1 on Wed Mar 22 20:50:28 2023
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO fullchip
  CLASS BLOCK ;
  SIZE 474.400000 BY 473.600000 ;
  FOREIGN fullchip 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 178.150000 0.600000 178.250000 ;
    END
  END clk
  PIN mem_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 294.150000 0.600000 294.250000 ;
    END
  END mem_in[127]
  PIN mem_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 293.350000 0.600000 293.450000 ;
    END
  END mem_in[126]
  PIN mem_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 292.550000 0.600000 292.650000 ;
    END
  END mem_in[125]
  PIN mem_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 291.750000 0.600000 291.850000 ;
    END
  END mem_in[124]
  PIN mem_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 290.950000 0.600000 291.050000 ;
    END
  END mem_in[123]
  PIN mem_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 290.150000 0.600000 290.250000 ;
    END
  END mem_in[122]
  PIN mem_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 289.350000 0.600000 289.450000 ;
    END
  END mem_in[121]
  PIN mem_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 288.550000 0.600000 288.650000 ;
    END
  END mem_in[120]
  PIN mem_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 287.750000 0.600000 287.850000 ;
    END
  END mem_in[119]
  PIN mem_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 286.950000 0.600000 287.050000 ;
    END
  END mem_in[118]
  PIN mem_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 286.150000 0.600000 286.250000 ;
    END
  END mem_in[117]
  PIN mem_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 285.350000 0.600000 285.450000 ;
    END
  END mem_in[116]
  PIN mem_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 284.550000 0.600000 284.650000 ;
    END
  END mem_in[115]
  PIN mem_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 283.750000 0.600000 283.850000 ;
    END
  END mem_in[114]
  PIN mem_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 282.950000 0.600000 283.050000 ;
    END
  END mem_in[113]
  PIN mem_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 282.150000 0.600000 282.250000 ;
    END
  END mem_in[112]
  PIN mem_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 281.350000 0.600000 281.450000 ;
    END
  END mem_in[111]
  PIN mem_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 280.550000 0.600000 280.650000 ;
    END
  END mem_in[110]
  PIN mem_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 279.750000 0.600000 279.850000 ;
    END
  END mem_in[109]
  PIN mem_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 278.950000 0.600000 279.050000 ;
    END
  END mem_in[108]
  PIN mem_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 278.150000 0.600000 278.250000 ;
    END
  END mem_in[107]
  PIN mem_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 277.350000 0.600000 277.450000 ;
    END
  END mem_in[106]
  PIN mem_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 276.550000 0.600000 276.650000 ;
    END
  END mem_in[105]
  PIN mem_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 275.750000 0.600000 275.850000 ;
    END
  END mem_in[104]
  PIN mem_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 274.950000 0.600000 275.050000 ;
    END
  END mem_in[103]
  PIN mem_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 274.150000 0.600000 274.250000 ;
    END
  END mem_in[102]
  PIN mem_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 273.350000 0.600000 273.450000 ;
    END
  END mem_in[101]
  PIN mem_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 272.550000 0.600000 272.650000 ;
    END
  END mem_in[100]
  PIN mem_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 271.750000 0.600000 271.850000 ;
    END
  END mem_in[99]
  PIN mem_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 270.950000 0.600000 271.050000 ;
    END
  END mem_in[98]
  PIN mem_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 270.150000 0.600000 270.250000 ;
    END
  END mem_in[97]
  PIN mem_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 269.350000 0.600000 269.450000 ;
    END
  END mem_in[96]
  PIN mem_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 268.550000 0.600000 268.650000 ;
    END
  END mem_in[95]
  PIN mem_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 267.750000 0.600000 267.850000 ;
    END
  END mem_in[94]
  PIN mem_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 266.950000 0.600000 267.050000 ;
    END
  END mem_in[93]
  PIN mem_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 266.150000 0.600000 266.250000 ;
    END
  END mem_in[92]
  PIN mem_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 265.350000 0.600000 265.450000 ;
    END
  END mem_in[91]
  PIN mem_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 264.550000 0.600000 264.650000 ;
    END
  END mem_in[90]
  PIN mem_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 263.750000 0.600000 263.850000 ;
    END
  END mem_in[89]
  PIN mem_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 262.950000 0.600000 263.050000 ;
    END
  END mem_in[88]
  PIN mem_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 262.150000 0.600000 262.250000 ;
    END
  END mem_in[87]
  PIN mem_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 261.350000 0.600000 261.450000 ;
    END
  END mem_in[86]
  PIN mem_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 260.550000 0.600000 260.650000 ;
    END
  END mem_in[85]
  PIN mem_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 259.750000 0.600000 259.850000 ;
    END
  END mem_in[84]
  PIN mem_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 258.950000 0.600000 259.050000 ;
    END
  END mem_in[83]
  PIN mem_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 258.150000 0.600000 258.250000 ;
    END
  END mem_in[82]
  PIN mem_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 257.350000 0.600000 257.450000 ;
    END
  END mem_in[81]
  PIN mem_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 256.550000 0.600000 256.650000 ;
    END
  END mem_in[80]
  PIN mem_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 255.750000 0.600000 255.850000 ;
    END
  END mem_in[79]
  PIN mem_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 254.950000 0.600000 255.050000 ;
    END
  END mem_in[78]
  PIN mem_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 254.150000 0.600000 254.250000 ;
    END
  END mem_in[77]
  PIN mem_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 253.350000 0.600000 253.450000 ;
    END
  END mem_in[76]
  PIN mem_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 252.550000 0.600000 252.650000 ;
    END
  END mem_in[75]
  PIN mem_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 251.750000 0.600000 251.850000 ;
    END
  END mem_in[74]
  PIN mem_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 250.950000 0.600000 251.050000 ;
    END
  END mem_in[73]
  PIN mem_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 250.150000 0.600000 250.250000 ;
    END
  END mem_in[72]
  PIN mem_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 249.350000 0.600000 249.450000 ;
    END
  END mem_in[71]
  PIN mem_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 248.550000 0.600000 248.650000 ;
    END
  END mem_in[70]
  PIN mem_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 247.750000 0.600000 247.850000 ;
    END
  END mem_in[69]
  PIN mem_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 246.950000 0.600000 247.050000 ;
    END
  END mem_in[68]
  PIN mem_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 246.150000 0.600000 246.250000 ;
    END
  END mem_in[67]
  PIN mem_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 245.350000 0.600000 245.450000 ;
    END
  END mem_in[66]
  PIN mem_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 244.550000 0.600000 244.650000 ;
    END
  END mem_in[65]
  PIN mem_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 243.750000 0.600000 243.850000 ;
    END
  END mem_in[64]
  PIN mem_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 242.950000 0.600000 243.050000 ;
    END
  END mem_in[63]
  PIN mem_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 242.150000 0.600000 242.250000 ;
    END
  END mem_in[62]
  PIN mem_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 241.350000 0.600000 241.450000 ;
    END
  END mem_in[61]
  PIN mem_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 240.550000 0.600000 240.650000 ;
    END
  END mem_in[60]
  PIN mem_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 239.750000 0.600000 239.850000 ;
    END
  END mem_in[59]
  PIN mem_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 238.950000 0.600000 239.050000 ;
    END
  END mem_in[58]
  PIN mem_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 238.150000 0.600000 238.250000 ;
    END
  END mem_in[57]
  PIN mem_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 237.350000 0.600000 237.450000 ;
    END
  END mem_in[56]
  PIN mem_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 236.550000 0.600000 236.650000 ;
    END
  END mem_in[55]
  PIN mem_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 235.750000 0.600000 235.850000 ;
    END
  END mem_in[54]
  PIN mem_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 234.950000 0.600000 235.050000 ;
    END
  END mem_in[53]
  PIN mem_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 234.150000 0.600000 234.250000 ;
    END
  END mem_in[52]
  PIN mem_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 233.350000 0.600000 233.450000 ;
    END
  END mem_in[51]
  PIN mem_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 232.550000 0.600000 232.650000 ;
    END
  END mem_in[50]
  PIN mem_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 231.750000 0.600000 231.850000 ;
    END
  END mem_in[49]
  PIN mem_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 230.950000 0.600000 231.050000 ;
    END
  END mem_in[48]
  PIN mem_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 230.150000 0.600000 230.250000 ;
    END
  END mem_in[47]
  PIN mem_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 229.350000 0.600000 229.450000 ;
    END
  END mem_in[46]
  PIN mem_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 228.550000 0.600000 228.650000 ;
    END
  END mem_in[45]
  PIN mem_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 227.750000 0.600000 227.850000 ;
    END
  END mem_in[44]
  PIN mem_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 226.950000 0.600000 227.050000 ;
    END
  END mem_in[43]
  PIN mem_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 226.150000 0.600000 226.250000 ;
    END
  END mem_in[42]
  PIN mem_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 225.350000 0.600000 225.450000 ;
    END
  END mem_in[41]
  PIN mem_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 224.550000 0.600000 224.650000 ;
    END
  END mem_in[40]
  PIN mem_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 223.750000 0.600000 223.850000 ;
    END
  END mem_in[39]
  PIN mem_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 222.950000 0.600000 223.050000 ;
    END
  END mem_in[38]
  PIN mem_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 222.150000 0.600000 222.250000 ;
    END
  END mem_in[37]
  PIN mem_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 221.350000 0.600000 221.450000 ;
    END
  END mem_in[36]
  PIN mem_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 220.550000 0.600000 220.650000 ;
    END
  END mem_in[35]
  PIN mem_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 219.750000 0.600000 219.850000 ;
    END
  END mem_in[34]
  PIN mem_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 218.950000 0.600000 219.050000 ;
    END
  END mem_in[33]
  PIN mem_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 218.150000 0.600000 218.250000 ;
    END
  END mem_in[32]
  PIN mem_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 217.350000 0.600000 217.450000 ;
    END
  END mem_in[31]
  PIN mem_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 216.550000 0.600000 216.650000 ;
    END
  END mem_in[30]
  PIN mem_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 215.750000 0.600000 215.850000 ;
    END
  END mem_in[29]
  PIN mem_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 214.950000 0.600000 215.050000 ;
    END
  END mem_in[28]
  PIN mem_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 214.150000 0.600000 214.250000 ;
    END
  END mem_in[27]
  PIN mem_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 213.350000 0.600000 213.450000 ;
    END
  END mem_in[26]
  PIN mem_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 212.550000 0.600000 212.650000 ;
    END
  END mem_in[25]
  PIN mem_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 211.750000 0.600000 211.850000 ;
    END
  END mem_in[24]
  PIN mem_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 210.950000 0.600000 211.050000 ;
    END
  END mem_in[23]
  PIN mem_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 210.150000 0.600000 210.250000 ;
    END
  END mem_in[22]
  PIN mem_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 209.350000 0.600000 209.450000 ;
    END
  END mem_in[21]
  PIN mem_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 208.550000 0.600000 208.650000 ;
    END
  END mem_in[20]
  PIN mem_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 207.750000 0.600000 207.850000 ;
    END
  END mem_in[19]
  PIN mem_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 206.950000 0.600000 207.050000 ;
    END
  END mem_in[18]
  PIN mem_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 206.150000 0.600000 206.250000 ;
    END
  END mem_in[17]
  PIN mem_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 205.350000 0.600000 205.450000 ;
    END
  END mem_in[16]
  PIN mem_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 204.550000 0.600000 204.650000 ;
    END
  END mem_in[15]
  PIN mem_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 203.750000 0.600000 203.850000 ;
    END
  END mem_in[14]
  PIN mem_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 202.950000 0.600000 203.050000 ;
    END
  END mem_in[13]
  PIN mem_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 202.150000 0.600000 202.250000 ;
    END
  END mem_in[12]
  PIN mem_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 201.350000 0.600000 201.450000 ;
    END
  END mem_in[11]
  PIN mem_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 200.550000 0.600000 200.650000 ;
    END
  END mem_in[10]
  PIN mem_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 199.750000 0.600000 199.850000 ;
    END
  END mem_in[9]
  PIN mem_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 198.950000 0.600000 199.050000 ;
    END
  END mem_in[8]
  PIN mem_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 198.150000 0.600000 198.250000 ;
    END
  END mem_in[7]
  PIN mem_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 197.350000 0.600000 197.450000 ;
    END
  END mem_in[6]
  PIN mem_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 196.550000 0.600000 196.650000 ;
    END
  END mem_in[5]
  PIN mem_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 195.750000 0.600000 195.850000 ;
    END
  END mem_in[4]
  PIN mem_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 194.950000 0.600000 195.050000 ;
    END
  END mem_in[3]
  PIN mem_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 194.150000 0.600000 194.250000 ;
    END
  END mem_in[2]
  PIN mem_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 193.350000 0.600000 193.450000 ;
    END
  END mem_in[1]
  PIN mem_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 192.550000 0.600000 192.650000 ;
    END
  END mem_in[0]
  PIN inst[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 191.750000 0.600000 191.850000 ;
    END
  END inst[16]
  PIN inst[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 190.950000 0.600000 191.050000 ;
    END
  END inst[15]
  PIN inst[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 190.150000 0.600000 190.250000 ;
    END
  END inst[14]
  PIN inst[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 189.350000 0.600000 189.450000 ;
    END
  END inst[13]
  PIN inst[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 188.550000 0.600000 188.650000 ;
    END
  END inst[12]
  PIN inst[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 187.750000 0.600000 187.850000 ;
    END
  END inst[11]
  PIN inst[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 186.950000 0.600000 187.050000 ;
    END
  END inst[10]
  PIN inst[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 186.150000 0.600000 186.250000 ;
    END
  END inst[9]
  PIN inst[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 185.350000 0.600000 185.450000 ;
    END
  END inst[8]
  PIN inst[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 184.550000 0.600000 184.650000 ;
    END
  END inst[7]
  PIN inst[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 183.750000 0.600000 183.850000 ;
    END
  END inst[6]
  PIN inst[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 182.950000 0.600000 183.050000 ;
    END
  END inst[5]
  PIN inst[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 182.150000 0.600000 182.250000 ;
    END
  END inst[4]
  PIN inst[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 181.350000 0.600000 181.450000 ;
    END
  END inst[3]
  PIN inst[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 180.550000 0.600000 180.650000 ;
    END
  END inst[2]
  PIN inst[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 179.750000 0.600000 179.850000 ;
    END
  END inst[1]
  PIN inst[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 178.950000 0.600000 179.050000 ;
    END
  END inst[0]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 294.950000 0.600000 295.050000 ;
    END
  END reset
  PIN out[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 173.350000 474.400000 173.450000 ;
    END
  END out[159]
  PIN out[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 174.150000 474.400000 174.250000 ;
    END
  END out[158]
  PIN out[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 174.950000 474.400000 175.050000 ;
    END
  END out[157]
  PIN out[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 175.750000 474.400000 175.850000 ;
    END
  END out[156]
  PIN out[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 176.550000 474.400000 176.650000 ;
    END
  END out[155]
  PIN out[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 177.350000 474.400000 177.450000 ;
    END
  END out[154]
  PIN out[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 178.150000 474.400000 178.250000 ;
    END
  END out[153]
  PIN out[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 178.950000 474.400000 179.050000 ;
    END
  END out[152]
  PIN out[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 179.750000 474.400000 179.850000 ;
    END
  END out[151]
  PIN out[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 180.550000 474.400000 180.650000 ;
    END
  END out[150]
  PIN out[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 181.350000 474.400000 181.450000 ;
    END
  END out[149]
  PIN out[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 182.150000 474.400000 182.250000 ;
    END
  END out[148]
  PIN out[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 182.950000 474.400000 183.050000 ;
    END
  END out[147]
  PIN out[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 183.750000 474.400000 183.850000 ;
    END
  END out[146]
  PIN out[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 184.550000 474.400000 184.650000 ;
    END
  END out[145]
  PIN out[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 185.350000 474.400000 185.450000 ;
    END
  END out[144]
  PIN out[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 186.150000 474.400000 186.250000 ;
    END
  END out[143]
  PIN out[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 186.950000 474.400000 187.050000 ;
    END
  END out[142]
  PIN out[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 187.750000 474.400000 187.850000 ;
    END
  END out[141]
  PIN out[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 188.550000 474.400000 188.650000 ;
    END
  END out[140]
  PIN out[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 189.350000 474.400000 189.450000 ;
    END
  END out[139]
  PIN out[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 190.150000 474.400000 190.250000 ;
    END
  END out[138]
  PIN out[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 190.950000 474.400000 191.050000 ;
    END
  END out[137]
  PIN out[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 191.750000 474.400000 191.850000 ;
    END
  END out[136]
  PIN out[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 192.550000 474.400000 192.650000 ;
    END
  END out[135]
  PIN out[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 193.350000 474.400000 193.450000 ;
    END
  END out[134]
  PIN out[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 194.150000 474.400000 194.250000 ;
    END
  END out[133]
  PIN out[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 194.950000 474.400000 195.050000 ;
    END
  END out[132]
  PIN out[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 195.750000 474.400000 195.850000 ;
    END
  END out[131]
  PIN out[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 196.550000 474.400000 196.650000 ;
    END
  END out[130]
  PIN out[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 197.350000 474.400000 197.450000 ;
    END
  END out[129]
  PIN out[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 198.150000 474.400000 198.250000 ;
    END
  END out[128]
  PIN out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 198.950000 474.400000 199.050000 ;
    END
  END out[127]
  PIN out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 199.750000 474.400000 199.850000 ;
    END
  END out[126]
  PIN out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 200.550000 474.400000 200.650000 ;
    END
  END out[125]
  PIN out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 201.350000 474.400000 201.450000 ;
    END
  END out[124]
  PIN out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 202.150000 474.400000 202.250000 ;
    END
  END out[123]
  PIN out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 202.950000 474.400000 203.050000 ;
    END
  END out[122]
  PIN out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 203.750000 474.400000 203.850000 ;
    END
  END out[121]
  PIN out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 204.550000 474.400000 204.650000 ;
    END
  END out[120]
  PIN out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 205.350000 474.400000 205.450000 ;
    END
  END out[119]
  PIN out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 206.150000 474.400000 206.250000 ;
    END
  END out[118]
  PIN out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 206.950000 474.400000 207.050000 ;
    END
  END out[117]
  PIN out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 207.750000 474.400000 207.850000 ;
    END
  END out[116]
  PIN out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 208.550000 474.400000 208.650000 ;
    END
  END out[115]
  PIN out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 209.350000 474.400000 209.450000 ;
    END
  END out[114]
  PIN out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 210.150000 474.400000 210.250000 ;
    END
  END out[113]
  PIN out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 210.950000 474.400000 211.050000 ;
    END
  END out[112]
  PIN out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 211.750000 474.400000 211.850000 ;
    END
  END out[111]
  PIN out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 212.550000 474.400000 212.650000 ;
    END
  END out[110]
  PIN out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 213.350000 474.400000 213.450000 ;
    END
  END out[109]
  PIN out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 214.150000 474.400000 214.250000 ;
    END
  END out[108]
  PIN out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 214.950000 474.400000 215.050000 ;
    END
  END out[107]
  PIN out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 215.750000 474.400000 215.850000 ;
    END
  END out[106]
  PIN out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 216.550000 474.400000 216.650000 ;
    END
  END out[105]
  PIN out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 217.350000 474.400000 217.450000 ;
    END
  END out[104]
  PIN out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 218.150000 474.400000 218.250000 ;
    END
  END out[103]
  PIN out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 218.950000 474.400000 219.050000 ;
    END
  END out[102]
  PIN out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 219.750000 474.400000 219.850000 ;
    END
  END out[101]
  PIN out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 220.550000 474.400000 220.650000 ;
    END
  END out[100]
  PIN out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 221.350000 474.400000 221.450000 ;
    END
  END out[99]
  PIN out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 222.150000 474.400000 222.250000 ;
    END
  END out[98]
  PIN out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 222.950000 474.400000 223.050000 ;
    END
  END out[97]
  PIN out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 223.750000 474.400000 223.850000 ;
    END
  END out[96]
  PIN out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 224.550000 474.400000 224.650000 ;
    END
  END out[95]
  PIN out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 225.350000 474.400000 225.450000 ;
    END
  END out[94]
  PIN out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 226.150000 474.400000 226.250000 ;
    END
  END out[93]
  PIN out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 226.950000 474.400000 227.050000 ;
    END
  END out[92]
  PIN out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 227.750000 474.400000 227.850000 ;
    END
  END out[91]
  PIN out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 228.550000 474.400000 228.650000 ;
    END
  END out[90]
  PIN out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 229.350000 474.400000 229.450000 ;
    END
  END out[89]
  PIN out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 230.150000 474.400000 230.250000 ;
    END
  END out[88]
  PIN out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 230.950000 474.400000 231.050000 ;
    END
  END out[87]
  PIN out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 231.750000 474.400000 231.850000 ;
    END
  END out[86]
  PIN out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 232.550000 474.400000 232.650000 ;
    END
  END out[85]
  PIN out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 233.350000 474.400000 233.450000 ;
    END
  END out[84]
  PIN out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 234.150000 474.400000 234.250000 ;
    END
  END out[83]
  PIN out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 234.950000 474.400000 235.050000 ;
    END
  END out[82]
  PIN out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 235.750000 474.400000 235.850000 ;
    END
  END out[81]
  PIN out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 236.550000 474.400000 236.650000 ;
    END
  END out[80]
  PIN out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 237.350000 474.400000 237.450000 ;
    END
  END out[79]
  PIN out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 238.150000 474.400000 238.250000 ;
    END
  END out[78]
  PIN out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 238.950000 474.400000 239.050000 ;
    END
  END out[77]
  PIN out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 239.750000 474.400000 239.850000 ;
    END
  END out[76]
  PIN out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 240.550000 474.400000 240.650000 ;
    END
  END out[75]
  PIN out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 241.350000 474.400000 241.450000 ;
    END
  END out[74]
  PIN out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 242.150000 474.400000 242.250000 ;
    END
  END out[73]
  PIN out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 242.950000 474.400000 243.050000 ;
    END
  END out[72]
  PIN out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 243.750000 474.400000 243.850000 ;
    END
  END out[71]
  PIN out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 244.550000 474.400000 244.650000 ;
    END
  END out[70]
  PIN out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 245.350000 474.400000 245.450000 ;
    END
  END out[69]
  PIN out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 246.150000 474.400000 246.250000 ;
    END
  END out[68]
  PIN out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 246.950000 474.400000 247.050000 ;
    END
  END out[67]
  PIN out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 247.750000 474.400000 247.850000 ;
    END
  END out[66]
  PIN out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 248.550000 474.400000 248.650000 ;
    END
  END out[65]
  PIN out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 249.350000 474.400000 249.450000 ;
    END
  END out[64]
  PIN out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 250.150000 474.400000 250.250000 ;
    END
  END out[63]
  PIN out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 250.950000 474.400000 251.050000 ;
    END
  END out[62]
  PIN out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 251.750000 474.400000 251.850000 ;
    END
  END out[61]
  PIN out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 252.550000 474.400000 252.650000 ;
    END
  END out[60]
  PIN out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 253.350000 474.400000 253.450000 ;
    END
  END out[59]
  PIN out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 254.150000 474.400000 254.250000 ;
    END
  END out[58]
  PIN out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 254.950000 474.400000 255.050000 ;
    END
  END out[57]
  PIN out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 255.750000 474.400000 255.850000 ;
    END
  END out[56]
  PIN out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 256.550000 474.400000 256.650000 ;
    END
  END out[55]
  PIN out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 257.350000 474.400000 257.450000 ;
    END
  END out[54]
  PIN out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 258.150000 474.400000 258.250000 ;
    END
  END out[53]
  PIN out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 258.950000 474.400000 259.050000 ;
    END
  END out[52]
  PIN out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 259.750000 474.400000 259.850000 ;
    END
  END out[51]
  PIN out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 260.550000 474.400000 260.650000 ;
    END
  END out[50]
  PIN out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 261.350000 474.400000 261.450000 ;
    END
  END out[49]
  PIN out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 262.150000 474.400000 262.250000 ;
    END
  END out[48]
  PIN out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 262.950000 474.400000 263.050000 ;
    END
  END out[47]
  PIN out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 263.750000 474.400000 263.850000 ;
    END
  END out[46]
  PIN out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 264.550000 474.400000 264.650000 ;
    END
  END out[45]
  PIN out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 265.350000 474.400000 265.450000 ;
    END
  END out[44]
  PIN out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 266.150000 474.400000 266.250000 ;
    END
  END out[43]
  PIN out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 266.950000 474.400000 267.050000 ;
    END
  END out[42]
  PIN out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 267.750000 474.400000 267.850000 ;
    END
  END out[41]
  PIN out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 268.550000 474.400000 268.650000 ;
    END
  END out[40]
  PIN out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 269.350000 474.400000 269.450000 ;
    END
  END out[39]
  PIN out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 270.150000 474.400000 270.250000 ;
    END
  END out[38]
  PIN out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 270.950000 474.400000 271.050000 ;
    END
  END out[37]
  PIN out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 271.750000 474.400000 271.850000 ;
    END
  END out[36]
  PIN out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 272.550000 474.400000 272.650000 ;
    END
  END out[35]
  PIN out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 273.350000 474.400000 273.450000 ;
    END
  END out[34]
  PIN out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 274.150000 474.400000 274.250000 ;
    END
  END out[33]
  PIN out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 274.950000 474.400000 275.050000 ;
    END
  END out[32]
  PIN out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 275.750000 474.400000 275.850000 ;
    END
  END out[31]
  PIN out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 276.550000 474.400000 276.650000 ;
    END
  END out[30]
  PIN out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 277.350000 474.400000 277.450000 ;
    END
  END out[29]
  PIN out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 278.150000 474.400000 278.250000 ;
    END
  END out[28]
  PIN out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 278.950000 474.400000 279.050000 ;
    END
  END out[27]
  PIN out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 279.750000 474.400000 279.850000 ;
    END
  END out[26]
  PIN out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 280.550000 474.400000 280.650000 ;
    END
  END out[25]
  PIN out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 281.350000 474.400000 281.450000 ;
    END
  END out[24]
  PIN out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 282.150000 474.400000 282.250000 ;
    END
  END out[23]
  PIN out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 282.950000 474.400000 283.050000 ;
    END
  END out[22]
  PIN out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 283.750000 474.400000 283.850000 ;
    END
  END out[21]
  PIN out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 284.550000 474.400000 284.650000 ;
    END
  END out[20]
  PIN out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 285.350000 474.400000 285.450000 ;
    END
  END out[19]
  PIN out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 286.150000 474.400000 286.250000 ;
    END
  END out[18]
  PIN out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 286.950000 474.400000 287.050000 ;
    END
  END out[17]
  PIN out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 287.750000 474.400000 287.850000 ;
    END
  END out[16]
  PIN out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 288.550000 474.400000 288.650000 ;
    END
  END out[15]
  PIN out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 289.350000 474.400000 289.450000 ;
    END
  END out[14]
  PIN out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 290.150000 474.400000 290.250000 ;
    END
  END out[13]
  PIN out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 290.950000 474.400000 291.050000 ;
    END
  END out[12]
  PIN out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 291.750000 474.400000 291.850000 ;
    END
  END out[11]
  PIN out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 292.550000 474.400000 292.650000 ;
    END
  END out[10]
  PIN out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 293.350000 474.400000 293.450000 ;
    END
  END out[9]
  PIN out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 294.150000 474.400000 294.250000 ;
    END
  END out[8]
  PIN out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 294.950000 474.400000 295.050000 ;
    END
  END out[7]
  PIN out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 295.750000 474.400000 295.850000 ;
    END
  END out[6]
  PIN out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 296.550000 474.400000 296.650000 ;
    END
  END out[5]
  PIN out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 297.350000 474.400000 297.450000 ;
    END
  END out[4]
  PIN out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 298.150000 474.400000 298.250000 ;
    END
  END out[3]
  PIN out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 298.950000 474.400000 299.050000 ;
    END
  END out[2]
  PIN out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 299.750000 474.400000 299.850000 ;
    END
  END out[1]
  PIN out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.800000 300.550000 474.400000 300.650000 ;
    END
  END out[0]
  OBS
    LAYER M1 ;
      RECT 0.000000 0.000000 474.400000 473.600000 ;
    LAYER M2 ;
      RECT 0.000000 0.000000 474.400000 473.600000 ;
    LAYER M3 ;
      RECT 0.000000 300.750000 474.400000 473.600000 ;
      RECT 0.000000 300.450000 473.680000 300.750000 ;
      RECT 0.000000 299.950000 474.400000 300.450000 ;
      RECT 0.000000 299.650000 473.680000 299.950000 ;
      RECT 0.000000 299.150000 474.400000 299.650000 ;
      RECT 0.000000 298.850000 473.680000 299.150000 ;
      RECT 0.000000 298.350000 474.400000 298.850000 ;
      RECT 0.000000 298.050000 473.680000 298.350000 ;
      RECT 0.000000 297.550000 474.400000 298.050000 ;
      RECT 0.000000 297.250000 473.680000 297.550000 ;
      RECT 0.000000 296.750000 474.400000 297.250000 ;
      RECT 0.000000 296.450000 473.680000 296.750000 ;
      RECT 0.000000 295.950000 474.400000 296.450000 ;
      RECT 0.000000 295.650000 473.680000 295.950000 ;
      RECT 0.000000 295.150000 474.400000 295.650000 ;
      RECT 0.720000 294.850000 473.680000 295.150000 ;
      RECT 0.000000 294.350000 474.400000 294.850000 ;
      RECT 0.720000 294.050000 473.680000 294.350000 ;
      RECT 0.000000 293.550000 474.400000 294.050000 ;
      RECT 0.720000 293.250000 473.680000 293.550000 ;
      RECT 0.000000 292.750000 474.400000 293.250000 ;
      RECT 0.720000 292.450000 473.680000 292.750000 ;
      RECT 0.000000 291.950000 474.400000 292.450000 ;
      RECT 0.720000 291.650000 473.680000 291.950000 ;
      RECT 0.000000 291.150000 474.400000 291.650000 ;
      RECT 0.720000 290.850000 473.680000 291.150000 ;
      RECT 0.000000 290.350000 474.400000 290.850000 ;
      RECT 0.720000 290.050000 473.680000 290.350000 ;
      RECT 0.000000 289.550000 474.400000 290.050000 ;
      RECT 0.720000 289.250000 473.680000 289.550000 ;
      RECT 0.000000 288.750000 474.400000 289.250000 ;
      RECT 0.720000 288.450000 473.680000 288.750000 ;
      RECT 0.000000 287.950000 474.400000 288.450000 ;
      RECT 0.720000 287.650000 473.680000 287.950000 ;
      RECT 0.000000 287.150000 474.400000 287.650000 ;
      RECT 0.720000 286.850000 473.680000 287.150000 ;
      RECT 0.000000 286.350000 474.400000 286.850000 ;
      RECT 0.720000 286.050000 473.680000 286.350000 ;
      RECT 0.000000 285.550000 474.400000 286.050000 ;
      RECT 0.720000 285.250000 473.680000 285.550000 ;
      RECT 0.000000 284.750000 474.400000 285.250000 ;
      RECT 0.720000 284.450000 473.680000 284.750000 ;
      RECT 0.000000 283.950000 474.400000 284.450000 ;
      RECT 0.720000 283.650000 473.680000 283.950000 ;
      RECT 0.000000 283.150000 474.400000 283.650000 ;
      RECT 0.720000 282.850000 473.680000 283.150000 ;
      RECT 0.000000 282.350000 474.400000 282.850000 ;
      RECT 0.720000 282.050000 473.680000 282.350000 ;
      RECT 0.000000 281.550000 474.400000 282.050000 ;
      RECT 0.720000 281.250000 473.680000 281.550000 ;
      RECT 0.000000 280.750000 474.400000 281.250000 ;
      RECT 0.720000 280.450000 473.680000 280.750000 ;
      RECT 0.000000 279.950000 474.400000 280.450000 ;
      RECT 0.720000 279.650000 473.680000 279.950000 ;
      RECT 0.000000 279.150000 474.400000 279.650000 ;
      RECT 0.720000 278.850000 473.680000 279.150000 ;
      RECT 0.000000 278.350000 474.400000 278.850000 ;
      RECT 0.720000 278.050000 473.680000 278.350000 ;
      RECT 0.000000 277.550000 474.400000 278.050000 ;
      RECT 0.720000 277.250000 473.680000 277.550000 ;
      RECT 0.000000 276.750000 474.400000 277.250000 ;
      RECT 0.720000 276.450000 473.680000 276.750000 ;
      RECT 0.000000 275.950000 474.400000 276.450000 ;
      RECT 0.720000 275.650000 473.680000 275.950000 ;
      RECT 0.000000 275.150000 474.400000 275.650000 ;
      RECT 0.720000 274.850000 473.680000 275.150000 ;
      RECT 0.000000 274.350000 474.400000 274.850000 ;
      RECT 0.720000 274.050000 473.680000 274.350000 ;
      RECT 0.000000 273.550000 474.400000 274.050000 ;
      RECT 0.720000 273.250000 473.680000 273.550000 ;
      RECT 0.000000 272.750000 474.400000 273.250000 ;
      RECT 0.720000 272.450000 473.680000 272.750000 ;
      RECT 0.000000 271.950000 474.400000 272.450000 ;
      RECT 0.720000 271.650000 473.680000 271.950000 ;
      RECT 0.000000 271.150000 474.400000 271.650000 ;
      RECT 0.720000 270.850000 473.680000 271.150000 ;
      RECT 0.000000 270.350000 474.400000 270.850000 ;
      RECT 0.720000 270.050000 473.680000 270.350000 ;
      RECT 0.000000 269.550000 474.400000 270.050000 ;
      RECT 0.720000 269.250000 473.680000 269.550000 ;
      RECT 0.000000 268.750000 474.400000 269.250000 ;
      RECT 0.720000 268.450000 473.680000 268.750000 ;
      RECT 0.000000 267.950000 474.400000 268.450000 ;
      RECT 0.720000 267.650000 473.680000 267.950000 ;
      RECT 0.000000 267.150000 474.400000 267.650000 ;
      RECT 0.720000 266.850000 473.680000 267.150000 ;
      RECT 0.000000 266.350000 474.400000 266.850000 ;
      RECT 0.720000 266.050000 473.680000 266.350000 ;
      RECT 0.000000 265.550000 474.400000 266.050000 ;
      RECT 0.720000 265.250000 473.680000 265.550000 ;
      RECT 0.000000 264.750000 474.400000 265.250000 ;
      RECT 0.720000 264.450000 473.680000 264.750000 ;
      RECT 0.000000 263.950000 474.400000 264.450000 ;
      RECT 0.720000 263.650000 473.680000 263.950000 ;
      RECT 0.000000 263.150000 474.400000 263.650000 ;
      RECT 0.720000 262.850000 473.680000 263.150000 ;
      RECT 0.000000 262.350000 474.400000 262.850000 ;
      RECT 0.720000 262.050000 473.680000 262.350000 ;
      RECT 0.000000 261.550000 474.400000 262.050000 ;
      RECT 0.720000 261.250000 473.680000 261.550000 ;
      RECT 0.000000 260.750000 474.400000 261.250000 ;
      RECT 0.720000 260.450000 473.680000 260.750000 ;
      RECT 0.000000 259.950000 474.400000 260.450000 ;
      RECT 0.720000 259.650000 473.680000 259.950000 ;
      RECT 0.000000 259.150000 474.400000 259.650000 ;
      RECT 0.720000 258.850000 473.680000 259.150000 ;
      RECT 0.000000 258.350000 474.400000 258.850000 ;
      RECT 0.720000 258.050000 473.680000 258.350000 ;
      RECT 0.000000 257.550000 474.400000 258.050000 ;
      RECT 0.720000 257.250000 473.680000 257.550000 ;
      RECT 0.000000 256.750000 474.400000 257.250000 ;
      RECT 0.720000 256.450000 473.680000 256.750000 ;
      RECT 0.000000 255.950000 474.400000 256.450000 ;
      RECT 0.720000 255.650000 473.680000 255.950000 ;
      RECT 0.000000 255.150000 474.400000 255.650000 ;
      RECT 0.720000 254.850000 473.680000 255.150000 ;
      RECT 0.000000 254.350000 474.400000 254.850000 ;
      RECT 0.720000 254.050000 473.680000 254.350000 ;
      RECT 0.000000 253.550000 474.400000 254.050000 ;
      RECT 0.720000 253.250000 473.680000 253.550000 ;
      RECT 0.000000 252.750000 474.400000 253.250000 ;
      RECT 0.720000 252.450000 473.680000 252.750000 ;
      RECT 0.000000 251.950000 474.400000 252.450000 ;
      RECT 0.720000 251.650000 473.680000 251.950000 ;
      RECT 0.000000 251.150000 474.400000 251.650000 ;
      RECT 0.720000 250.850000 473.680000 251.150000 ;
      RECT 0.000000 250.350000 474.400000 250.850000 ;
      RECT 0.720000 250.050000 473.680000 250.350000 ;
      RECT 0.000000 249.550000 474.400000 250.050000 ;
      RECT 0.720000 249.250000 473.680000 249.550000 ;
      RECT 0.000000 248.750000 474.400000 249.250000 ;
      RECT 0.720000 248.450000 473.680000 248.750000 ;
      RECT 0.000000 247.950000 474.400000 248.450000 ;
      RECT 0.720000 247.650000 473.680000 247.950000 ;
      RECT 0.000000 247.150000 474.400000 247.650000 ;
      RECT 0.720000 246.850000 473.680000 247.150000 ;
      RECT 0.000000 246.350000 474.400000 246.850000 ;
      RECT 0.720000 246.050000 473.680000 246.350000 ;
      RECT 0.000000 245.550000 474.400000 246.050000 ;
      RECT 0.720000 245.250000 473.680000 245.550000 ;
      RECT 0.000000 244.750000 474.400000 245.250000 ;
      RECT 0.720000 244.450000 473.680000 244.750000 ;
      RECT 0.000000 243.950000 474.400000 244.450000 ;
      RECT 0.720000 243.650000 473.680000 243.950000 ;
      RECT 0.000000 243.150000 474.400000 243.650000 ;
      RECT 0.720000 242.850000 473.680000 243.150000 ;
      RECT 0.000000 242.350000 474.400000 242.850000 ;
      RECT 0.720000 242.050000 473.680000 242.350000 ;
      RECT 0.000000 241.550000 474.400000 242.050000 ;
      RECT 0.720000 241.250000 473.680000 241.550000 ;
      RECT 0.000000 240.750000 474.400000 241.250000 ;
      RECT 0.720000 240.450000 473.680000 240.750000 ;
      RECT 0.000000 239.950000 474.400000 240.450000 ;
      RECT 0.720000 239.650000 473.680000 239.950000 ;
      RECT 0.000000 239.150000 474.400000 239.650000 ;
      RECT 0.720000 238.850000 473.680000 239.150000 ;
      RECT 0.000000 238.350000 474.400000 238.850000 ;
      RECT 0.720000 238.050000 473.680000 238.350000 ;
      RECT 0.000000 237.550000 474.400000 238.050000 ;
      RECT 0.720000 237.250000 473.680000 237.550000 ;
      RECT 0.000000 236.750000 474.400000 237.250000 ;
      RECT 0.720000 236.450000 473.680000 236.750000 ;
      RECT 0.000000 235.950000 474.400000 236.450000 ;
      RECT 0.720000 235.650000 473.680000 235.950000 ;
      RECT 0.000000 235.150000 474.400000 235.650000 ;
      RECT 0.720000 234.850000 473.680000 235.150000 ;
      RECT 0.000000 234.350000 474.400000 234.850000 ;
      RECT 0.720000 234.050000 473.680000 234.350000 ;
      RECT 0.000000 233.550000 474.400000 234.050000 ;
      RECT 0.720000 233.250000 473.680000 233.550000 ;
      RECT 0.000000 232.750000 474.400000 233.250000 ;
      RECT 0.720000 232.450000 473.680000 232.750000 ;
      RECT 0.000000 231.950000 474.400000 232.450000 ;
      RECT 0.720000 231.650000 473.680000 231.950000 ;
      RECT 0.000000 231.150000 474.400000 231.650000 ;
      RECT 0.720000 230.850000 473.680000 231.150000 ;
      RECT 0.000000 230.350000 474.400000 230.850000 ;
      RECT 0.720000 230.050000 473.680000 230.350000 ;
      RECT 0.000000 229.550000 474.400000 230.050000 ;
      RECT 0.720000 229.250000 473.680000 229.550000 ;
      RECT 0.000000 228.750000 474.400000 229.250000 ;
      RECT 0.720000 228.450000 473.680000 228.750000 ;
      RECT 0.000000 227.950000 474.400000 228.450000 ;
      RECT 0.720000 227.650000 473.680000 227.950000 ;
      RECT 0.000000 227.150000 474.400000 227.650000 ;
      RECT 0.720000 226.850000 473.680000 227.150000 ;
      RECT 0.000000 226.350000 474.400000 226.850000 ;
      RECT 0.720000 226.050000 473.680000 226.350000 ;
      RECT 0.000000 225.550000 474.400000 226.050000 ;
      RECT 0.720000 225.250000 473.680000 225.550000 ;
      RECT 0.000000 224.750000 474.400000 225.250000 ;
      RECT 0.720000 224.450000 473.680000 224.750000 ;
      RECT 0.000000 223.950000 474.400000 224.450000 ;
      RECT 0.720000 223.650000 473.680000 223.950000 ;
      RECT 0.000000 223.150000 474.400000 223.650000 ;
      RECT 0.720000 222.850000 473.680000 223.150000 ;
      RECT 0.000000 222.350000 474.400000 222.850000 ;
      RECT 0.720000 222.050000 473.680000 222.350000 ;
      RECT 0.000000 221.550000 474.400000 222.050000 ;
      RECT 0.720000 221.250000 473.680000 221.550000 ;
      RECT 0.000000 220.750000 474.400000 221.250000 ;
      RECT 0.720000 220.450000 473.680000 220.750000 ;
      RECT 0.000000 219.950000 474.400000 220.450000 ;
      RECT 0.720000 219.650000 473.680000 219.950000 ;
      RECT 0.000000 219.150000 474.400000 219.650000 ;
      RECT 0.720000 218.850000 473.680000 219.150000 ;
      RECT 0.000000 218.350000 474.400000 218.850000 ;
      RECT 0.720000 218.050000 473.680000 218.350000 ;
      RECT 0.000000 217.550000 474.400000 218.050000 ;
      RECT 0.720000 217.250000 473.680000 217.550000 ;
      RECT 0.000000 216.750000 474.400000 217.250000 ;
      RECT 0.720000 216.450000 473.680000 216.750000 ;
      RECT 0.000000 215.950000 474.400000 216.450000 ;
      RECT 0.720000 215.650000 473.680000 215.950000 ;
      RECT 0.000000 215.150000 474.400000 215.650000 ;
      RECT 0.720000 214.850000 473.680000 215.150000 ;
      RECT 0.000000 214.350000 474.400000 214.850000 ;
      RECT 0.720000 214.050000 473.680000 214.350000 ;
      RECT 0.000000 213.550000 474.400000 214.050000 ;
      RECT 0.720000 213.250000 473.680000 213.550000 ;
      RECT 0.000000 212.750000 474.400000 213.250000 ;
      RECT 0.720000 212.450000 473.680000 212.750000 ;
      RECT 0.000000 211.950000 474.400000 212.450000 ;
      RECT 0.720000 211.650000 473.680000 211.950000 ;
      RECT 0.000000 211.150000 474.400000 211.650000 ;
      RECT 0.720000 210.850000 473.680000 211.150000 ;
      RECT 0.000000 210.350000 474.400000 210.850000 ;
      RECT 0.720000 210.050000 473.680000 210.350000 ;
      RECT 0.000000 209.550000 474.400000 210.050000 ;
      RECT 0.720000 209.250000 473.680000 209.550000 ;
      RECT 0.000000 208.750000 474.400000 209.250000 ;
      RECT 0.720000 208.450000 473.680000 208.750000 ;
      RECT 0.000000 207.950000 474.400000 208.450000 ;
      RECT 0.720000 207.650000 473.680000 207.950000 ;
      RECT 0.000000 207.150000 474.400000 207.650000 ;
      RECT 0.720000 206.850000 473.680000 207.150000 ;
      RECT 0.000000 206.350000 474.400000 206.850000 ;
      RECT 0.720000 206.050000 473.680000 206.350000 ;
      RECT 0.000000 205.550000 474.400000 206.050000 ;
      RECT 0.720000 205.250000 473.680000 205.550000 ;
      RECT 0.000000 204.750000 474.400000 205.250000 ;
      RECT 0.720000 204.450000 473.680000 204.750000 ;
      RECT 0.000000 203.950000 474.400000 204.450000 ;
      RECT 0.720000 203.650000 473.680000 203.950000 ;
      RECT 0.000000 203.150000 474.400000 203.650000 ;
      RECT 0.720000 202.850000 473.680000 203.150000 ;
      RECT 0.000000 202.350000 474.400000 202.850000 ;
      RECT 0.720000 202.050000 473.680000 202.350000 ;
      RECT 0.000000 201.550000 474.400000 202.050000 ;
      RECT 0.720000 201.250000 473.680000 201.550000 ;
      RECT 0.000000 200.750000 474.400000 201.250000 ;
      RECT 0.720000 200.450000 473.680000 200.750000 ;
      RECT 0.000000 199.950000 474.400000 200.450000 ;
      RECT 0.720000 199.650000 473.680000 199.950000 ;
      RECT 0.000000 199.150000 474.400000 199.650000 ;
      RECT 0.720000 198.850000 473.680000 199.150000 ;
      RECT 0.000000 198.350000 474.400000 198.850000 ;
      RECT 0.720000 198.050000 473.680000 198.350000 ;
      RECT 0.000000 197.550000 474.400000 198.050000 ;
      RECT 0.720000 197.250000 473.680000 197.550000 ;
      RECT 0.000000 196.750000 474.400000 197.250000 ;
      RECT 0.720000 196.450000 473.680000 196.750000 ;
      RECT 0.000000 195.950000 474.400000 196.450000 ;
      RECT 0.720000 195.650000 473.680000 195.950000 ;
      RECT 0.000000 195.150000 474.400000 195.650000 ;
      RECT 0.720000 194.850000 473.680000 195.150000 ;
      RECT 0.000000 194.350000 474.400000 194.850000 ;
      RECT 0.720000 194.050000 473.680000 194.350000 ;
      RECT 0.000000 193.550000 474.400000 194.050000 ;
      RECT 0.720000 193.250000 473.680000 193.550000 ;
      RECT 0.000000 192.750000 474.400000 193.250000 ;
      RECT 0.720000 192.450000 473.680000 192.750000 ;
      RECT 0.000000 191.950000 474.400000 192.450000 ;
      RECT 0.720000 191.650000 473.680000 191.950000 ;
      RECT 0.000000 191.150000 474.400000 191.650000 ;
      RECT 0.720000 190.850000 473.680000 191.150000 ;
      RECT 0.000000 190.350000 474.400000 190.850000 ;
      RECT 0.720000 190.050000 473.680000 190.350000 ;
      RECT 0.000000 189.550000 474.400000 190.050000 ;
      RECT 0.720000 189.250000 473.680000 189.550000 ;
      RECT 0.000000 188.750000 474.400000 189.250000 ;
      RECT 0.720000 188.450000 473.680000 188.750000 ;
      RECT 0.000000 187.950000 474.400000 188.450000 ;
      RECT 0.720000 187.650000 473.680000 187.950000 ;
      RECT 0.000000 187.150000 474.400000 187.650000 ;
      RECT 0.720000 186.850000 473.680000 187.150000 ;
      RECT 0.000000 186.350000 474.400000 186.850000 ;
      RECT 0.720000 186.050000 473.680000 186.350000 ;
      RECT 0.000000 185.550000 474.400000 186.050000 ;
      RECT 0.720000 185.250000 473.680000 185.550000 ;
      RECT 0.000000 184.750000 474.400000 185.250000 ;
      RECT 0.720000 184.450000 473.680000 184.750000 ;
      RECT 0.000000 183.950000 474.400000 184.450000 ;
      RECT 0.720000 183.650000 473.680000 183.950000 ;
      RECT 0.000000 183.150000 474.400000 183.650000 ;
      RECT 0.720000 182.850000 473.680000 183.150000 ;
      RECT 0.000000 182.350000 474.400000 182.850000 ;
      RECT 0.720000 182.050000 473.680000 182.350000 ;
      RECT 0.000000 181.550000 474.400000 182.050000 ;
      RECT 0.720000 181.250000 473.680000 181.550000 ;
      RECT 0.000000 180.750000 474.400000 181.250000 ;
      RECT 0.720000 180.450000 473.680000 180.750000 ;
      RECT 0.000000 179.950000 474.400000 180.450000 ;
      RECT 0.720000 179.650000 473.680000 179.950000 ;
      RECT 0.000000 179.150000 474.400000 179.650000 ;
      RECT 0.720000 178.850000 473.680000 179.150000 ;
      RECT 0.000000 178.350000 474.400000 178.850000 ;
      RECT 0.720000 178.050000 473.680000 178.350000 ;
      RECT 0.000000 177.550000 474.400000 178.050000 ;
      RECT 0.000000 177.250000 473.680000 177.550000 ;
      RECT 0.000000 176.750000 474.400000 177.250000 ;
      RECT 0.000000 176.450000 473.680000 176.750000 ;
      RECT 0.000000 175.950000 474.400000 176.450000 ;
      RECT 0.000000 175.650000 473.680000 175.950000 ;
      RECT 0.000000 175.150000 474.400000 175.650000 ;
      RECT 0.000000 174.850000 473.680000 175.150000 ;
      RECT 0.000000 174.350000 474.400000 174.850000 ;
      RECT 0.000000 174.050000 473.680000 174.350000 ;
      RECT 0.000000 173.550000 474.400000 174.050000 ;
      RECT 0.000000 173.250000 473.680000 173.550000 ;
      RECT 0.000000 0.000000 474.400000 173.250000 ;
    LAYER M4 ;
      RECT 0.000000 0.000000 474.400000 473.600000 ;
    LAYER M5 ;
      RECT 0.000000 0.000000 474.400000 473.600000 ;
    LAYER M6 ;
      RECT 0.000000 0.000000 474.400000 473.600000 ;
    LAYER M7 ;
      RECT 0.000000 0.000000 474.400000 473.600000 ;
    LAYER M8 ;
      RECT 0.000000 0.000000 474.400000 473.600000 ;
  END
END fullchip

END LIBRARY
