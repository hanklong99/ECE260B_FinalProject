##
## LEF for PtnCells ;
## created by Innovus v19.17-s077_1 on Fri Mar 17 15:44:05 2023
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO fullchip
  CLASS BLOCK ;
  SIZE 679.200000 BY 677.000000 ;
  FOREIGN fullchip 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 263.550000 0.600000 263.650000 ;
    END
  END clk0
  PIN clk1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 264.350000 0.600000 264.450000 ;
    END
  END clk1
  PIN mem_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 411.550000 0.600000 411.650000 ;
    END
  END mem_in[63]
  PIN mem_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 410.750000 0.600000 410.850000 ;
    END
  END mem_in[62]
  PIN mem_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 409.950000 0.600000 410.050000 ;
    END
  END mem_in[61]
  PIN mem_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 409.150000 0.600000 409.250000 ;
    END
  END mem_in[60]
  PIN mem_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 408.350000 0.600000 408.450000 ;
    END
  END mem_in[59]
  PIN mem_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 407.550000 0.600000 407.650000 ;
    END
  END mem_in[58]
  PIN mem_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 406.750000 0.600000 406.850000 ;
    END
  END mem_in[57]
  PIN mem_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 405.950000 0.600000 406.050000 ;
    END
  END mem_in[56]
  PIN mem_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 405.150000 0.600000 405.250000 ;
    END
  END mem_in[55]
  PIN mem_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 404.350000 0.600000 404.450000 ;
    END
  END mem_in[54]
  PIN mem_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 403.550000 0.600000 403.650000 ;
    END
  END mem_in[53]
  PIN mem_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 402.750000 0.600000 402.850000 ;
    END
  END mem_in[52]
  PIN mem_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 401.950000 0.600000 402.050000 ;
    END
  END mem_in[51]
  PIN mem_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 401.150000 0.600000 401.250000 ;
    END
  END mem_in[50]
  PIN mem_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 400.350000 0.600000 400.450000 ;
    END
  END mem_in[49]
  PIN mem_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 399.550000 0.600000 399.650000 ;
    END
  END mem_in[48]
  PIN mem_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 398.750000 0.600000 398.850000 ;
    END
  END mem_in[47]
  PIN mem_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 397.950000 0.600000 398.050000 ;
    END
  END mem_in[46]
  PIN mem_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 397.150000 0.600000 397.250000 ;
    END
  END mem_in[45]
  PIN mem_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 396.350000 0.600000 396.450000 ;
    END
  END mem_in[44]
  PIN mem_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 395.550000 0.600000 395.650000 ;
    END
  END mem_in[43]
  PIN mem_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 394.750000 0.600000 394.850000 ;
    END
  END mem_in[42]
  PIN mem_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 393.950000 0.600000 394.050000 ;
    END
  END mem_in[41]
  PIN mem_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 393.150000 0.600000 393.250000 ;
    END
  END mem_in[40]
  PIN mem_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 392.350000 0.600000 392.450000 ;
    END
  END mem_in[39]
  PIN mem_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 391.550000 0.600000 391.650000 ;
    END
  END mem_in[38]
  PIN mem_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 390.750000 0.600000 390.850000 ;
    END
  END mem_in[37]
  PIN mem_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 389.950000 0.600000 390.050000 ;
    END
  END mem_in[36]
  PIN mem_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 389.150000 0.600000 389.250000 ;
    END
  END mem_in[35]
  PIN mem_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 388.350000 0.600000 388.450000 ;
    END
  END mem_in[34]
  PIN mem_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 387.550000 0.600000 387.650000 ;
    END
  END mem_in[33]
  PIN mem_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 386.750000 0.600000 386.850000 ;
    END
  END mem_in[32]
  PIN mem_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 385.950000 0.600000 386.050000 ;
    END
  END mem_in[31]
  PIN mem_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 385.150000 0.600000 385.250000 ;
    END
  END mem_in[30]
  PIN mem_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 384.350000 0.600000 384.450000 ;
    END
  END mem_in[29]
  PIN mem_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 383.550000 0.600000 383.650000 ;
    END
  END mem_in[28]
  PIN mem_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 382.750000 0.600000 382.850000 ;
    END
  END mem_in[27]
  PIN mem_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 381.950000 0.600000 382.050000 ;
    END
  END mem_in[26]
  PIN mem_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 381.150000 0.600000 381.250000 ;
    END
  END mem_in[25]
  PIN mem_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 380.350000 0.600000 380.450000 ;
    END
  END mem_in[24]
  PIN mem_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 379.550000 0.600000 379.650000 ;
    END
  END mem_in[23]
  PIN mem_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 378.750000 0.600000 378.850000 ;
    END
  END mem_in[22]
  PIN mem_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 377.950000 0.600000 378.050000 ;
    END
  END mem_in[21]
  PIN mem_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 377.150000 0.600000 377.250000 ;
    END
  END mem_in[20]
  PIN mem_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 376.350000 0.600000 376.450000 ;
    END
  END mem_in[19]
  PIN mem_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 375.550000 0.600000 375.650000 ;
    END
  END mem_in[18]
  PIN mem_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 374.750000 0.600000 374.850000 ;
    END
  END mem_in[17]
  PIN mem_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 373.950000 0.600000 374.050000 ;
    END
  END mem_in[16]
  PIN mem_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 373.150000 0.600000 373.250000 ;
    END
  END mem_in[15]
  PIN mem_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 372.350000 0.600000 372.450000 ;
    END
  END mem_in[14]
  PIN mem_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 371.550000 0.600000 371.650000 ;
    END
  END mem_in[13]
  PIN mem_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 370.750000 0.600000 370.850000 ;
    END
  END mem_in[12]
  PIN mem_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 369.950000 0.600000 370.050000 ;
    END
  END mem_in[11]
  PIN mem_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 369.150000 0.600000 369.250000 ;
    END
  END mem_in[10]
  PIN mem_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 368.350000 0.600000 368.450000 ;
    END
  END mem_in[9]
  PIN mem_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 367.550000 0.600000 367.650000 ;
    END
  END mem_in[8]
  PIN mem_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 366.750000 0.600000 366.850000 ;
    END
  END mem_in[7]
  PIN mem_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 365.950000 0.600000 366.050000 ;
    END
  END mem_in[6]
  PIN mem_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 365.150000 0.600000 365.250000 ;
    END
  END mem_in[5]
  PIN mem_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 364.350000 0.600000 364.450000 ;
    END
  END mem_in[4]
  PIN mem_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 363.550000 0.600000 363.650000 ;
    END
  END mem_in[3]
  PIN mem_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 362.750000 0.600000 362.850000 ;
    END
  END mem_in[2]
  PIN mem_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 361.950000 0.600000 362.050000 ;
    END
  END mem_in[1]
  PIN mem_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 361.150000 0.600000 361.250000 ;
    END
  END mem_in[0]
  PIN mem_in1[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 360.350000 0.600000 360.450000 ;
    END
  END mem_in1[63]
  PIN mem_in1[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 359.550000 0.600000 359.650000 ;
    END
  END mem_in1[62]
  PIN mem_in1[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 358.750000 0.600000 358.850000 ;
    END
  END mem_in1[61]
  PIN mem_in1[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 357.950000 0.600000 358.050000 ;
    END
  END mem_in1[60]
  PIN mem_in1[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 357.150000 0.600000 357.250000 ;
    END
  END mem_in1[59]
  PIN mem_in1[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 356.350000 0.600000 356.450000 ;
    END
  END mem_in1[58]
  PIN mem_in1[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 355.550000 0.600000 355.650000 ;
    END
  END mem_in1[57]
  PIN mem_in1[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 354.750000 0.600000 354.850000 ;
    END
  END mem_in1[56]
  PIN mem_in1[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 353.950000 0.600000 354.050000 ;
    END
  END mem_in1[55]
  PIN mem_in1[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 353.150000 0.600000 353.250000 ;
    END
  END mem_in1[54]
  PIN mem_in1[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 352.350000 0.600000 352.450000 ;
    END
  END mem_in1[53]
  PIN mem_in1[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 351.550000 0.600000 351.650000 ;
    END
  END mem_in1[52]
  PIN mem_in1[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 350.750000 0.600000 350.850000 ;
    END
  END mem_in1[51]
  PIN mem_in1[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 349.950000 0.600000 350.050000 ;
    END
  END mem_in1[50]
  PIN mem_in1[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 349.150000 0.600000 349.250000 ;
    END
  END mem_in1[49]
  PIN mem_in1[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 348.350000 0.600000 348.450000 ;
    END
  END mem_in1[48]
  PIN mem_in1[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 347.550000 0.600000 347.650000 ;
    END
  END mem_in1[47]
  PIN mem_in1[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 346.750000 0.600000 346.850000 ;
    END
  END mem_in1[46]
  PIN mem_in1[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 345.950000 0.600000 346.050000 ;
    END
  END mem_in1[45]
  PIN mem_in1[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 345.150000 0.600000 345.250000 ;
    END
  END mem_in1[44]
  PIN mem_in1[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 344.350000 0.600000 344.450000 ;
    END
  END mem_in1[43]
  PIN mem_in1[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 343.550000 0.600000 343.650000 ;
    END
  END mem_in1[42]
  PIN mem_in1[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 342.750000 0.600000 342.850000 ;
    END
  END mem_in1[41]
  PIN mem_in1[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 341.950000 0.600000 342.050000 ;
    END
  END mem_in1[40]
  PIN mem_in1[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 341.150000 0.600000 341.250000 ;
    END
  END mem_in1[39]
  PIN mem_in1[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 340.350000 0.600000 340.450000 ;
    END
  END mem_in1[38]
  PIN mem_in1[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 339.550000 0.600000 339.650000 ;
    END
  END mem_in1[37]
  PIN mem_in1[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 338.750000 0.600000 338.850000 ;
    END
  END mem_in1[36]
  PIN mem_in1[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 337.950000 0.600000 338.050000 ;
    END
  END mem_in1[35]
  PIN mem_in1[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 337.150000 0.600000 337.250000 ;
    END
  END mem_in1[34]
  PIN mem_in1[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 336.350000 0.600000 336.450000 ;
    END
  END mem_in1[33]
  PIN mem_in1[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 335.550000 0.600000 335.650000 ;
    END
  END mem_in1[32]
  PIN mem_in1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 334.750000 0.600000 334.850000 ;
    END
  END mem_in1[31]
  PIN mem_in1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 333.950000 0.600000 334.050000 ;
    END
  END mem_in1[30]
  PIN mem_in1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 333.150000 0.600000 333.250000 ;
    END
  END mem_in1[29]
  PIN mem_in1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 332.350000 0.600000 332.450000 ;
    END
  END mem_in1[28]
  PIN mem_in1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 331.550000 0.600000 331.650000 ;
    END
  END mem_in1[27]
  PIN mem_in1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 330.750000 0.600000 330.850000 ;
    END
  END mem_in1[26]
  PIN mem_in1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 329.950000 0.600000 330.050000 ;
    END
  END mem_in1[25]
  PIN mem_in1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 329.150000 0.600000 329.250000 ;
    END
  END mem_in1[24]
  PIN mem_in1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 328.350000 0.600000 328.450000 ;
    END
  END mem_in1[23]
  PIN mem_in1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 327.550000 0.600000 327.650000 ;
    END
  END mem_in1[22]
  PIN mem_in1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 326.750000 0.600000 326.850000 ;
    END
  END mem_in1[21]
  PIN mem_in1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 325.950000 0.600000 326.050000 ;
    END
  END mem_in1[20]
  PIN mem_in1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 325.150000 0.600000 325.250000 ;
    END
  END mem_in1[19]
  PIN mem_in1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 324.350000 0.600000 324.450000 ;
    END
  END mem_in1[18]
  PIN mem_in1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 323.550000 0.600000 323.650000 ;
    END
  END mem_in1[17]
  PIN mem_in1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 322.750000 0.600000 322.850000 ;
    END
  END mem_in1[16]
  PIN mem_in1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 321.950000 0.600000 322.050000 ;
    END
  END mem_in1[15]
  PIN mem_in1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 321.150000 0.600000 321.250000 ;
    END
  END mem_in1[14]
  PIN mem_in1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 320.350000 0.600000 320.450000 ;
    END
  END mem_in1[13]
  PIN mem_in1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 319.550000 0.600000 319.650000 ;
    END
  END mem_in1[12]
  PIN mem_in1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 318.750000 0.600000 318.850000 ;
    END
  END mem_in1[11]
  PIN mem_in1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 317.950000 0.600000 318.050000 ;
    END
  END mem_in1[10]
  PIN mem_in1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 317.150000 0.600000 317.250000 ;
    END
  END mem_in1[9]
  PIN mem_in1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 316.350000 0.600000 316.450000 ;
    END
  END mem_in1[8]
  PIN mem_in1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 315.550000 0.600000 315.650000 ;
    END
  END mem_in1[7]
  PIN mem_in1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 314.750000 0.600000 314.850000 ;
    END
  END mem_in1[6]
  PIN mem_in1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 313.950000 0.600000 314.050000 ;
    END
  END mem_in1[5]
  PIN mem_in1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 313.150000 0.600000 313.250000 ;
    END
  END mem_in1[4]
  PIN mem_in1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 312.350000 0.600000 312.450000 ;
    END
  END mem_in1[3]
  PIN mem_in1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 311.550000 0.600000 311.650000 ;
    END
  END mem_in1[2]
  PIN mem_in1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 310.750000 0.600000 310.850000 ;
    END
  END mem_in1[1]
  PIN mem_in1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 309.950000 0.600000 310.050000 ;
    END
  END mem_in1[0]
  PIN inst[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 309.150000 0.600000 309.250000 ;
    END
  END inst[27]
  PIN inst[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 308.350000 0.600000 308.450000 ;
    END
  END inst[26]
  PIN inst[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 307.550000 0.600000 307.650000 ;
    END
  END inst[25]
  PIN inst[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 306.750000 0.600000 306.850000 ;
    END
  END inst[24]
  PIN inst[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 305.950000 0.600000 306.050000 ;
    END
  END inst[23]
  PIN inst[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 305.150000 0.600000 305.250000 ;
    END
  END inst[22]
  PIN inst[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 304.350000 0.600000 304.450000 ;
    END
  END inst[21]
  PIN inst[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 303.550000 0.600000 303.650000 ;
    END
  END inst[20]
  PIN inst[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 302.750000 0.600000 302.850000 ;
    END
  END inst[19]
  PIN inst[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 301.950000 0.600000 302.050000 ;
    END
  END inst[18]
  PIN inst[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 301.150000 0.600000 301.250000 ;
    END
  END inst[17]
  PIN inst[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 300.350000 0.600000 300.450000 ;
    END
  END inst[16]
  PIN inst[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 299.550000 0.600000 299.650000 ;
    END
  END inst[15]
  PIN inst[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 298.750000 0.600000 298.850000 ;
    END
  END inst[14]
  PIN inst[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 297.950000 0.600000 298.050000 ;
    END
  END inst[13]
  PIN inst[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 297.150000 0.600000 297.250000 ;
    END
  END inst[12]
  PIN inst[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 296.350000 0.600000 296.450000 ;
    END
  END inst[11]
  PIN inst[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 295.550000 0.600000 295.650000 ;
    END
  END inst[10]
  PIN inst[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 294.750000 0.600000 294.850000 ;
    END
  END inst[9]
  PIN inst[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 293.950000 0.600000 294.050000 ;
    END
  END inst[8]
  PIN inst[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 293.150000 0.600000 293.250000 ;
    END
  END inst[7]
  PIN inst[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 292.350000 0.600000 292.450000 ;
    END
  END inst[6]
  PIN inst[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 291.550000 0.600000 291.650000 ;
    END
  END inst[5]
  PIN inst[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 290.750000 0.600000 290.850000 ;
    END
  END inst[4]
  PIN inst[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 289.950000 0.600000 290.050000 ;
    END
  END inst[3]
  PIN inst[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 289.150000 0.600000 289.250000 ;
    END
  END inst[2]
  PIN inst[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 288.350000 0.600000 288.450000 ;
    END
  END inst[1]
  PIN inst[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 287.550000 0.600000 287.650000 ;
    END
  END inst[0]
  PIN inst1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 286.750000 0.600000 286.850000 ;
    END
  END inst1[27]
  PIN inst1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 285.950000 0.600000 286.050000 ;
    END
  END inst1[26]
  PIN inst1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 285.150000 0.600000 285.250000 ;
    END
  END inst1[25]
  PIN inst1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 284.350000 0.600000 284.450000 ;
    END
  END inst1[24]
  PIN inst1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 283.550000 0.600000 283.650000 ;
    END
  END inst1[23]
  PIN inst1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 282.750000 0.600000 282.850000 ;
    END
  END inst1[22]
  PIN inst1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 281.950000 0.600000 282.050000 ;
    END
  END inst1[21]
  PIN inst1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 281.150000 0.600000 281.250000 ;
    END
  END inst1[20]
  PIN inst1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 280.350000 0.600000 280.450000 ;
    END
  END inst1[19]
  PIN inst1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 279.550000 0.600000 279.650000 ;
    END
  END inst1[18]
  PIN inst1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 278.750000 0.600000 278.850000 ;
    END
  END inst1[17]
  PIN inst1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 277.950000 0.600000 278.050000 ;
    END
  END inst1[16]
  PIN inst1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 277.150000 0.600000 277.250000 ;
    END
  END inst1[15]
  PIN inst1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 276.350000 0.600000 276.450000 ;
    END
  END inst1[14]
  PIN inst1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 275.550000 0.600000 275.650000 ;
    END
  END inst1[13]
  PIN inst1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 274.750000 0.600000 274.850000 ;
    END
  END inst1[12]
  PIN inst1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 273.950000 0.600000 274.050000 ;
    END
  END inst1[11]
  PIN inst1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 273.150000 0.600000 273.250000 ;
    END
  END inst1[10]
  PIN inst1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 272.350000 0.600000 272.450000 ;
    END
  END inst1[9]
  PIN inst1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 271.550000 0.600000 271.650000 ;
    END
  END inst1[8]
  PIN inst1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 270.750000 0.600000 270.850000 ;
    END
  END inst1[7]
  PIN inst1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 269.950000 0.600000 270.050000 ;
    END
  END inst1[6]
  PIN inst1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 269.150000 0.600000 269.250000 ;
    END
  END inst1[5]
  PIN inst1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 268.350000 0.600000 268.450000 ;
    END
  END inst1[4]
  PIN inst1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 267.550000 0.600000 267.650000 ;
    END
  END inst1[3]
  PIN inst1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 266.750000 0.600000 266.850000 ;
    END
  END inst1[2]
  PIN inst1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 265.950000 0.600000 266.050000 ;
    END
  END inst1[1]
  PIN inst1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 265.150000 0.600000 265.250000 ;
    END
  END inst1[0]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 412.350000 0.600000 412.450000 ;
    END
  END reset
  PIN reset1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 413.150000 0.600000 413.250000 ;
    END
  END reset1
  PIN out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 390.250000 0.000000 390.350000 0.600000 ;
    END
  END out[127]
  PIN out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 389.450000 0.000000 389.550000 0.600000 ;
    END
  END out[126]
  PIN out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 388.650000 0.000000 388.750000 0.600000 ;
    END
  END out[125]
  PIN out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 387.850000 0.000000 387.950000 0.600000 ;
    END
  END out[124]
  PIN out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 387.050000 0.000000 387.150000 0.600000 ;
    END
  END out[123]
  PIN out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 386.250000 0.000000 386.350000 0.600000 ;
    END
  END out[122]
  PIN out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 385.450000 0.000000 385.550000 0.600000 ;
    END
  END out[121]
  PIN out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 384.650000 0.000000 384.750000 0.600000 ;
    END
  END out[120]
  PIN out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 383.850000 0.000000 383.950000 0.600000 ;
    END
  END out[119]
  PIN out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 383.050000 0.000000 383.150000 0.600000 ;
    END
  END out[118]
  PIN out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.250000 0.000000 382.350000 0.600000 ;
    END
  END out[117]
  PIN out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 381.450000 0.000000 381.550000 0.600000 ;
    END
  END out[116]
  PIN out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 380.650000 0.000000 380.750000 0.600000 ;
    END
  END out[115]
  PIN out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 379.850000 0.000000 379.950000 0.600000 ;
    END
  END out[114]
  PIN out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 379.050000 0.000000 379.150000 0.600000 ;
    END
  END out[113]
  PIN out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 378.250000 0.000000 378.350000 0.600000 ;
    END
  END out[112]
  PIN out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 377.450000 0.000000 377.550000 0.600000 ;
    END
  END out[111]
  PIN out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 376.650000 0.000000 376.750000 0.600000 ;
    END
  END out[110]
  PIN out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 375.850000 0.000000 375.950000 0.600000 ;
    END
  END out[109]
  PIN out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 375.050000 0.000000 375.150000 0.600000 ;
    END
  END out[108]
  PIN out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 374.250000 0.000000 374.350000 0.600000 ;
    END
  END out[107]
  PIN out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 373.450000 0.000000 373.550000 0.600000 ;
    END
  END out[106]
  PIN out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 372.650000 0.000000 372.750000 0.600000 ;
    END
  END out[105]
  PIN out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 371.850000 0.000000 371.950000 0.600000 ;
    END
  END out[104]
  PIN out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 371.050000 0.000000 371.150000 0.600000 ;
    END
  END out[103]
  PIN out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 370.250000 0.000000 370.350000 0.600000 ;
    END
  END out[102]
  PIN out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 369.450000 0.000000 369.550000 0.600000 ;
    END
  END out[101]
  PIN out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 368.650000 0.000000 368.750000 0.600000 ;
    END
  END out[100]
  PIN out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 367.850000 0.000000 367.950000 0.600000 ;
    END
  END out[99]
  PIN out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 367.050000 0.000000 367.150000 0.600000 ;
    END
  END out[98]
  PIN out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 366.250000 0.000000 366.350000 0.600000 ;
    END
  END out[97]
  PIN out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 365.450000 0.000000 365.550000 0.600000 ;
    END
  END out[96]
  PIN out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 364.650000 0.000000 364.750000 0.600000 ;
    END
  END out[95]
  PIN out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 363.850000 0.000000 363.950000 0.600000 ;
    END
  END out[94]
  PIN out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 363.050000 0.000000 363.150000 0.600000 ;
    END
  END out[93]
  PIN out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 362.250000 0.000000 362.350000 0.600000 ;
    END
  END out[92]
  PIN out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 361.450000 0.000000 361.550000 0.600000 ;
    END
  END out[91]
  PIN out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 360.650000 0.000000 360.750000 0.600000 ;
    END
  END out[90]
  PIN out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 359.850000 0.000000 359.950000 0.600000 ;
    END
  END out[89]
  PIN out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 359.050000 0.000000 359.150000 0.600000 ;
    END
  END out[88]
  PIN out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 358.250000 0.000000 358.350000 0.600000 ;
    END
  END out[87]
  PIN out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 357.450000 0.000000 357.550000 0.600000 ;
    END
  END out[86]
  PIN out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 356.650000 0.000000 356.750000 0.600000 ;
    END
  END out[85]
  PIN out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 355.850000 0.000000 355.950000 0.600000 ;
    END
  END out[84]
  PIN out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 355.050000 0.000000 355.150000 0.600000 ;
    END
  END out[83]
  PIN out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 354.250000 0.000000 354.350000 0.600000 ;
    END
  END out[82]
  PIN out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 353.450000 0.000000 353.550000 0.600000 ;
    END
  END out[81]
  PIN out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 352.650000 0.000000 352.750000 0.600000 ;
    END
  END out[80]
  PIN out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 351.850000 0.000000 351.950000 0.600000 ;
    END
  END out[79]
  PIN out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 351.050000 0.000000 351.150000 0.600000 ;
    END
  END out[78]
  PIN out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 350.250000 0.000000 350.350000 0.600000 ;
    END
  END out[77]
  PIN out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 349.450000 0.000000 349.550000 0.600000 ;
    END
  END out[76]
  PIN out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 348.650000 0.000000 348.750000 0.600000 ;
    END
  END out[75]
  PIN out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 347.850000 0.000000 347.950000 0.600000 ;
    END
  END out[74]
  PIN out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 347.050000 0.000000 347.150000 0.600000 ;
    END
  END out[73]
  PIN out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 346.250000 0.000000 346.350000 0.600000 ;
    END
  END out[72]
  PIN out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 345.450000 0.000000 345.550000 0.600000 ;
    END
  END out[71]
  PIN out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 344.650000 0.000000 344.750000 0.600000 ;
    END
  END out[70]
  PIN out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 343.850000 0.000000 343.950000 0.600000 ;
    END
  END out[69]
  PIN out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 343.050000 0.000000 343.150000 0.600000 ;
    END
  END out[68]
  PIN out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 342.250000 0.000000 342.350000 0.600000 ;
    END
  END out[67]
  PIN out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 341.450000 0.000000 341.550000 0.600000 ;
    END
  END out[66]
  PIN out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 340.650000 0.000000 340.750000 0.600000 ;
    END
  END out[65]
  PIN out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 339.850000 0.000000 339.950000 0.600000 ;
    END
  END out[64]
  PIN out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 339.050000 0.000000 339.150000 0.600000 ;
    END
  END out[63]
  PIN out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 338.250000 0.000000 338.350000 0.600000 ;
    END
  END out[62]
  PIN out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 337.450000 0.000000 337.550000 0.600000 ;
    END
  END out[61]
  PIN out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 336.650000 0.000000 336.750000 0.600000 ;
    END
  END out[60]
  PIN out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 335.850000 0.000000 335.950000 0.600000 ;
    END
  END out[59]
  PIN out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 335.050000 0.000000 335.150000 0.600000 ;
    END
  END out[58]
  PIN out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 334.250000 0.000000 334.350000 0.600000 ;
    END
  END out[57]
  PIN out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 333.450000 0.000000 333.550000 0.600000 ;
    END
  END out[56]
  PIN out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 332.650000 0.000000 332.750000 0.600000 ;
    END
  END out[55]
  PIN out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 331.850000 0.000000 331.950000 0.600000 ;
    END
  END out[54]
  PIN out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 331.050000 0.000000 331.150000 0.600000 ;
    END
  END out[53]
  PIN out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 330.250000 0.000000 330.350000 0.600000 ;
    END
  END out[52]
  PIN out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 329.450000 0.000000 329.550000 0.600000 ;
    END
  END out[51]
  PIN out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 328.650000 0.000000 328.750000 0.600000 ;
    END
  END out[50]
  PIN out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 327.850000 0.000000 327.950000 0.600000 ;
    END
  END out[49]
  PIN out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 327.050000 0.000000 327.150000 0.600000 ;
    END
  END out[48]
  PIN out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 326.250000 0.000000 326.350000 0.600000 ;
    END
  END out[47]
  PIN out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 325.450000 0.000000 325.550000 0.600000 ;
    END
  END out[46]
  PIN out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 324.650000 0.000000 324.750000 0.600000 ;
    END
  END out[45]
  PIN out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 323.850000 0.000000 323.950000 0.600000 ;
    END
  END out[44]
  PIN out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 323.050000 0.000000 323.150000 0.600000 ;
    END
  END out[43]
  PIN out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 322.250000 0.000000 322.350000 0.600000 ;
    END
  END out[42]
  PIN out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 321.450000 0.000000 321.550000 0.600000 ;
    END
  END out[41]
  PIN out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 320.650000 0.000000 320.750000 0.600000 ;
    END
  END out[40]
  PIN out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 319.850000 0.000000 319.950000 0.600000 ;
    END
  END out[39]
  PIN out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 319.050000 0.000000 319.150000 0.600000 ;
    END
  END out[38]
  PIN out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 318.250000 0.000000 318.350000 0.600000 ;
    END
  END out[37]
  PIN out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 317.450000 0.000000 317.550000 0.600000 ;
    END
  END out[36]
  PIN out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 316.650000 0.000000 316.750000 0.600000 ;
    END
  END out[35]
  PIN out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 315.850000 0.000000 315.950000 0.600000 ;
    END
  END out[34]
  PIN out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 315.050000 0.000000 315.150000 0.600000 ;
    END
  END out[33]
  PIN out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 314.250000 0.000000 314.350000 0.600000 ;
    END
  END out[32]
  PIN out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 313.450000 0.000000 313.550000 0.600000 ;
    END
  END out[31]
  PIN out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 312.650000 0.000000 312.750000 0.600000 ;
    END
  END out[30]
  PIN out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 311.850000 0.000000 311.950000 0.600000 ;
    END
  END out[29]
  PIN out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 311.050000 0.000000 311.150000 0.600000 ;
    END
  END out[28]
  PIN out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 310.250000 0.000000 310.350000 0.600000 ;
    END
  END out[27]
  PIN out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 309.450000 0.000000 309.550000 0.600000 ;
    END
  END out[26]
  PIN out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 308.650000 0.000000 308.750000 0.600000 ;
    END
  END out[25]
  PIN out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 307.850000 0.000000 307.950000 0.600000 ;
    END
  END out[24]
  PIN out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 307.050000 0.000000 307.150000 0.600000 ;
    END
  END out[23]
  PIN out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 306.250000 0.000000 306.350000 0.600000 ;
    END
  END out[22]
  PIN out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 305.450000 0.000000 305.550000 0.600000 ;
    END
  END out[21]
  PIN out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 304.650000 0.000000 304.750000 0.600000 ;
    END
  END out[20]
  PIN out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 303.850000 0.000000 303.950000 0.600000 ;
    END
  END out[19]
  PIN out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 303.050000 0.000000 303.150000 0.600000 ;
    END
  END out[18]
  PIN out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 302.250000 0.000000 302.350000 0.600000 ;
    END
  END out[17]
  PIN out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 301.450000 0.000000 301.550000 0.600000 ;
    END
  END out[16]
  PIN out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 300.650000 0.000000 300.750000 0.600000 ;
    END
  END out[15]
  PIN out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 299.850000 0.000000 299.950000 0.600000 ;
    END
  END out[14]
  PIN out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 299.050000 0.000000 299.150000 0.600000 ;
    END
  END out[13]
  PIN out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 298.250000 0.000000 298.350000 0.600000 ;
    END
  END out[12]
  PIN out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 297.450000 0.000000 297.550000 0.600000 ;
    END
  END out[11]
  PIN out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 296.650000 0.000000 296.750000 0.600000 ;
    END
  END out[10]
  PIN out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 295.850000 0.000000 295.950000 0.600000 ;
    END
  END out[9]
  PIN out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 295.050000 0.000000 295.150000 0.600000 ;
    END
  END out[8]
  PIN out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 294.250000 0.000000 294.350000 0.600000 ;
    END
  END out[7]
  PIN out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 293.450000 0.000000 293.550000 0.600000 ;
    END
  END out[6]
  PIN out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 292.650000 0.000000 292.750000 0.600000 ;
    END
  END out[5]
  PIN out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 291.850000 0.000000 291.950000 0.600000 ;
    END
  END out[4]
  PIN out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 291.050000 0.000000 291.150000 0.600000 ;
    END
  END out[3]
  PIN out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 290.250000 0.000000 290.350000 0.600000 ;
    END
  END out[2]
  PIN out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 289.450000 0.000000 289.550000 0.600000 ;
    END
  END out[1]
  PIN out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 288.650000 0.000000 288.750000 0.600000 ;
    END
  END out[0]
  OBS
    LAYER M1 ;
      RECT 0.000000 0.000000 679.200000 677.000000 ;
    LAYER M2 ;
      RECT 0.000000 0.000000 679.200000 677.000000 ;
    LAYER M3 ;
      RECT 0.000000 413.350000 679.200000 677.000000 ;
      RECT 0.720000 413.050000 679.200000 413.350000 ;
      RECT 0.000000 412.550000 679.200000 413.050000 ;
      RECT 0.720000 412.250000 679.200000 412.550000 ;
      RECT 0.000000 411.750000 679.200000 412.250000 ;
      RECT 0.720000 411.450000 679.200000 411.750000 ;
      RECT 0.000000 410.950000 679.200000 411.450000 ;
      RECT 0.720000 410.650000 679.200000 410.950000 ;
      RECT 0.000000 410.150000 679.200000 410.650000 ;
      RECT 0.720000 409.850000 679.200000 410.150000 ;
      RECT 0.000000 409.350000 679.200000 409.850000 ;
      RECT 0.720000 409.050000 679.200000 409.350000 ;
      RECT 0.000000 408.550000 679.200000 409.050000 ;
      RECT 0.720000 408.250000 679.200000 408.550000 ;
      RECT 0.000000 407.750000 679.200000 408.250000 ;
      RECT 0.720000 407.450000 679.200000 407.750000 ;
      RECT 0.000000 406.950000 679.200000 407.450000 ;
      RECT 0.720000 406.650000 679.200000 406.950000 ;
      RECT 0.000000 406.150000 679.200000 406.650000 ;
      RECT 0.720000 405.850000 679.200000 406.150000 ;
      RECT 0.000000 405.350000 679.200000 405.850000 ;
      RECT 0.720000 405.050000 679.200000 405.350000 ;
      RECT 0.000000 404.550000 679.200000 405.050000 ;
      RECT 0.720000 404.250000 679.200000 404.550000 ;
      RECT 0.000000 403.750000 679.200000 404.250000 ;
      RECT 0.720000 403.450000 679.200000 403.750000 ;
      RECT 0.000000 402.950000 679.200000 403.450000 ;
      RECT 0.720000 402.650000 679.200000 402.950000 ;
      RECT 0.000000 402.150000 679.200000 402.650000 ;
      RECT 0.720000 401.850000 679.200000 402.150000 ;
      RECT 0.000000 401.350000 679.200000 401.850000 ;
      RECT 0.720000 401.050000 679.200000 401.350000 ;
      RECT 0.000000 400.550000 679.200000 401.050000 ;
      RECT 0.720000 400.250000 679.200000 400.550000 ;
      RECT 0.000000 399.750000 679.200000 400.250000 ;
      RECT 0.720000 399.450000 679.200000 399.750000 ;
      RECT 0.000000 398.950000 679.200000 399.450000 ;
      RECT 0.720000 398.650000 679.200000 398.950000 ;
      RECT 0.000000 398.150000 679.200000 398.650000 ;
      RECT 0.720000 397.850000 679.200000 398.150000 ;
      RECT 0.000000 397.350000 679.200000 397.850000 ;
      RECT 0.720000 397.050000 679.200000 397.350000 ;
      RECT 0.000000 396.550000 679.200000 397.050000 ;
      RECT 0.720000 396.250000 679.200000 396.550000 ;
      RECT 0.000000 395.750000 679.200000 396.250000 ;
      RECT 0.720000 395.450000 679.200000 395.750000 ;
      RECT 0.000000 394.950000 679.200000 395.450000 ;
      RECT 0.720000 394.650000 679.200000 394.950000 ;
      RECT 0.000000 394.150000 679.200000 394.650000 ;
      RECT 0.720000 393.850000 679.200000 394.150000 ;
      RECT 0.000000 393.350000 679.200000 393.850000 ;
      RECT 0.720000 393.050000 679.200000 393.350000 ;
      RECT 0.000000 392.550000 679.200000 393.050000 ;
      RECT 0.720000 392.250000 679.200000 392.550000 ;
      RECT 0.000000 391.750000 679.200000 392.250000 ;
      RECT 0.720000 391.450000 679.200000 391.750000 ;
      RECT 0.000000 390.950000 679.200000 391.450000 ;
      RECT 0.720000 390.650000 679.200000 390.950000 ;
      RECT 0.000000 390.150000 679.200000 390.650000 ;
      RECT 0.720000 389.850000 679.200000 390.150000 ;
      RECT 0.000000 389.350000 679.200000 389.850000 ;
      RECT 0.720000 389.050000 679.200000 389.350000 ;
      RECT 0.000000 388.550000 679.200000 389.050000 ;
      RECT 0.720000 388.250000 679.200000 388.550000 ;
      RECT 0.000000 387.750000 679.200000 388.250000 ;
      RECT 0.720000 387.450000 679.200000 387.750000 ;
      RECT 0.000000 386.950000 679.200000 387.450000 ;
      RECT 0.720000 386.650000 679.200000 386.950000 ;
      RECT 0.000000 386.150000 679.200000 386.650000 ;
      RECT 0.720000 385.850000 679.200000 386.150000 ;
      RECT 0.000000 385.350000 679.200000 385.850000 ;
      RECT 0.720000 385.050000 679.200000 385.350000 ;
      RECT 0.000000 384.550000 679.200000 385.050000 ;
      RECT 0.720000 384.250000 679.200000 384.550000 ;
      RECT 0.000000 383.750000 679.200000 384.250000 ;
      RECT 0.720000 383.450000 679.200000 383.750000 ;
      RECT 0.000000 382.950000 679.200000 383.450000 ;
      RECT 0.720000 382.650000 679.200000 382.950000 ;
      RECT 0.000000 382.150000 679.200000 382.650000 ;
      RECT 0.720000 381.850000 679.200000 382.150000 ;
      RECT 0.000000 381.350000 679.200000 381.850000 ;
      RECT 0.720000 381.050000 679.200000 381.350000 ;
      RECT 0.000000 380.550000 679.200000 381.050000 ;
      RECT 0.720000 380.250000 679.200000 380.550000 ;
      RECT 0.000000 379.750000 679.200000 380.250000 ;
      RECT 0.720000 379.450000 679.200000 379.750000 ;
      RECT 0.000000 378.950000 679.200000 379.450000 ;
      RECT 0.720000 378.650000 679.200000 378.950000 ;
      RECT 0.000000 378.150000 679.200000 378.650000 ;
      RECT 0.720000 377.850000 679.200000 378.150000 ;
      RECT 0.000000 377.350000 679.200000 377.850000 ;
      RECT 0.720000 377.050000 679.200000 377.350000 ;
      RECT 0.000000 376.550000 679.200000 377.050000 ;
      RECT 0.720000 376.250000 679.200000 376.550000 ;
      RECT 0.000000 375.750000 679.200000 376.250000 ;
      RECT 0.720000 375.450000 679.200000 375.750000 ;
      RECT 0.000000 374.950000 679.200000 375.450000 ;
      RECT 0.720000 374.650000 679.200000 374.950000 ;
      RECT 0.000000 374.150000 679.200000 374.650000 ;
      RECT 0.720000 373.850000 679.200000 374.150000 ;
      RECT 0.000000 373.350000 679.200000 373.850000 ;
      RECT 0.720000 373.050000 679.200000 373.350000 ;
      RECT 0.000000 372.550000 679.200000 373.050000 ;
      RECT 0.720000 372.250000 679.200000 372.550000 ;
      RECT 0.000000 371.750000 679.200000 372.250000 ;
      RECT 0.720000 371.450000 679.200000 371.750000 ;
      RECT 0.000000 370.950000 679.200000 371.450000 ;
      RECT 0.720000 370.650000 679.200000 370.950000 ;
      RECT 0.000000 370.150000 679.200000 370.650000 ;
      RECT 0.720000 369.850000 679.200000 370.150000 ;
      RECT 0.000000 369.350000 679.200000 369.850000 ;
      RECT 0.720000 369.050000 679.200000 369.350000 ;
      RECT 0.000000 368.550000 679.200000 369.050000 ;
      RECT 0.720000 368.250000 679.200000 368.550000 ;
      RECT 0.000000 367.750000 679.200000 368.250000 ;
      RECT 0.720000 367.450000 679.200000 367.750000 ;
      RECT 0.000000 366.950000 679.200000 367.450000 ;
      RECT 0.720000 366.650000 679.200000 366.950000 ;
      RECT 0.000000 366.150000 679.200000 366.650000 ;
      RECT 0.720000 365.850000 679.200000 366.150000 ;
      RECT 0.000000 365.350000 679.200000 365.850000 ;
      RECT 0.720000 365.050000 679.200000 365.350000 ;
      RECT 0.000000 364.550000 679.200000 365.050000 ;
      RECT 0.720000 364.250000 679.200000 364.550000 ;
      RECT 0.000000 363.750000 679.200000 364.250000 ;
      RECT 0.720000 363.450000 679.200000 363.750000 ;
      RECT 0.000000 362.950000 679.200000 363.450000 ;
      RECT 0.720000 362.650000 679.200000 362.950000 ;
      RECT 0.000000 362.150000 679.200000 362.650000 ;
      RECT 0.720000 361.850000 679.200000 362.150000 ;
      RECT 0.000000 361.350000 679.200000 361.850000 ;
      RECT 0.720000 361.050000 679.200000 361.350000 ;
      RECT 0.000000 360.550000 679.200000 361.050000 ;
      RECT 0.720000 360.250000 679.200000 360.550000 ;
      RECT 0.000000 359.750000 679.200000 360.250000 ;
      RECT 0.720000 359.450000 679.200000 359.750000 ;
      RECT 0.000000 358.950000 679.200000 359.450000 ;
      RECT 0.720000 358.650000 679.200000 358.950000 ;
      RECT 0.000000 358.150000 679.200000 358.650000 ;
      RECT 0.720000 357.850000 679.200000 358.150000 ;
      RECT 0.000000 357.350000 679.200000 357.850000 ;
      RECT 0.720000 357.050000 679.200000 357.350000 ;
      RECT 0.000000 356.550000 679.200000 357.050000 ;
      RECT 0.720000 356.250000 679.200000 356.550000 ;
      RECT 0.000000 355.750000 679.200000 356.250000 ;
      RECT 0.720000 355.450000 679.200000 355.750000 ;
      RECT 0.000000 354.950000 679.200000 355.450000 ;
      RECT 0.720000 354.650000 679.200000 354.950000 ;
      RECT 0.000000 354.150000 679.200000 354.650000 ;
      RECT 0.720000 353.850000 679.200000 354.150000 ;
      RECT 0.000000 353.350000 679.200000 353.850000 ;
      RECT 0.720000 353.050000 679.200000 353.350000 ;
      RECT 0.000000 352.550000 679.200000 353.050000 ;
      RECT 0.720000 352.250000 679.200000 352.550000 ;
      RECT 0.000000 351.750000 679.200000 352.250000 ;
      RECT 0.720000 351.450000 679.200000 351.750000 ;
      RECT 0.000000 350.950000 679.200000 351.450000 ;
      RECT 0.720000 350.650000 679.200000 350.950000 ;
      RECT 0.000000 350.150000 679.200000 350.650000 ;
      RECT 0.720000 349.850000 679.200000 350.150000 ;
      RECT 0.000000 349.350000 679.200000 349.850000 ;
      RECT 0.720000 349.050000 679.200000 349.350000 ;
      RECT 0.000000 348.550000 679.200000 349.050000 ;
      RECT 0.720000 348.250000 679.200000 348.550000 ;
      RECT 0.000000 347.750000 679.200000 348.250000 ;
      RECT 0.720000 347.450000 679.200000 347.750000 ;
      RECT 0.000000 346.950000 679.200000 347.450000 ;
      RECT 0.720000 346.650000 679.200000 346.950000 ;
      RECT 0.000000 346.150000 679.200000 346.650000 ;
      RECT 0.720000 345.850000 679.200000 346.150000 ;
      RECT 0.000000 345.350000 679.200000 345.850000 ;
      RECT 0.720000 345.050000 679.200000 345.350000 ;
      RECT 0.000000 344.550000 679.200000 345.050000 ;
      RECT 0.720000 344.250000 679.200000 344.550000 ;
      RECT 0.000000 343.750000 679.200000 344.250000 ;
      RECT 0.720000 343.450000 679.200000 343.750000 ;
      RECT 0.000000 342.950000 679.200000 343.450000 ;
      RECT 0.720000 342.650000 679.200000 342.950000 ;
      RECT 0.000000 342.150000 679.200000 342.650000 ;
      RECT 0.720000 341.850000 679.200000 342.150000 ;
      RECT 0.000000 341.350000 679.200000 341.850000 ;
      RECT 0.720000 341.050000 679.200000 341.350000 ;
      RECT 0.000000 340.550000 679.200000 341.050000 ;
      RECT 0.720000 340.250000 679.200000 340.550000 ;
      RECT 0.000000 339.750000 679.200000 340.250000 ;
      RECT 0.720000 339.450000 679.200000 339.750000 ;
      RECT 0.000000 338.950000 679.200000 339.450000 ;
      RECT 0.720000 338.650000 679.200000 338.950000 ;
      RECT 0.000000 338.150000 679.200000 338.650000 ;
      RECT 0.720000 337.850000 679.200000 338.150000 ;
      RECT 0.000000 337.350000 679.200000 337.850000 ;
      RECT 0.720000 337.050000 679.200000 337.350000 ;
      RECT 0.000000 336.550000 679.200000 337.050000 ;
      RECT 0.720000 336.250000 679.200000 336.550000 ;
      RECT 0.000000 335.750000 679.200000 336.250000 ;
      RECT 0.720000 335.450000 679.200000 335.750000 ;
      RECT 0.000000 334.950000 679.200000 335.450000 ;
      RECT 0.720000 334.650000 679.200000 334.950000 ;
      RECT 0.000000 334.150000 679.200000 334.650000 ;
      RECT 0.720000 333.850000 679.200000 334.150000 ;
      RECT 0.000000 333.350000 679.200000 333.850000 ;
      RECT 0.720000 333.050000 679.200000 333.350000 ;
      RECT 0.000000 332.550000 679.200000 333.050000 ;
      RECT 0.720000 332.250000 679.200000 332.550000 ;
      RECT 0.000000 331.750000 679.200000 332.250000 ;
      RECT 0.720000 331.450000 679.200000 331.750000 ;
      RECT 0.000000 330.950000 679.200000 331.450000 ;
      RECT 0.720000 330.650000 679.200000 330.950000 ;
      RECT 0.000000 330.150000 679.200000 330.650000 ;
      RECT 0.720000 329.850000 679.200000 330.150000 ;
      RECT 0.000000 329.350000 679.200000 329.850000 ;
      RECT 0.720000 329.050000 679.200000 329.350000 ;
      RECT 0.000000 328.550000 679.200000 329.050000 ;
      RECT 0.720000 328.250000 679.200000 328.550000 ;
      RECT 0.000000 327.750000 679.200000 328.250000 ;
      RECT 0.720000 327.450000 679.200000 327.750000 ;
      RECT 0.000000 326.950000 679.200000 327.450000 ;
      RECT 0.720000 326.650000 679.200000 326.950000 ;
      RECT 0.000000 326.150000 679.200000 326.650000 ;
      RECT 0.720000 325.850000 679.200000 326.150000 ;
      RECT 0.000000 325.350000 679.200000 325.850000 ;
      RECT 0.720000 325.050000 679.200000 325.350000 ;
      RECT 0.000000 324.550000 679.200000 325.050000 ;
      RECT 0.720000 324.250000 679.200000 324.550000 ;
      RECT 0.000000 323.750000 679.200000 324.250000 ;
      RECT 0.720000 323.450000 679.200000 323.750000 ;
      RECT 0.000000 322.950000 679.200000 323.450000 ;
      RECT 0.720000 322.650000 679.200000 322.950000 ;
      RECT 0.000000 322.150000 679.200000 322.650000 ;
      RECT 0.720000 321.850000 679.200000 322.150000 ;
      RECT 0.000000 321.350000 679.200000 321.850000 ;
      RECT 0.720000 321.050000 679.200000 321.350000 ;
      RECT 0.000000 320.550000 679.200000 321.050000 ;
      RECT 0.720000 320.250000 679.200000 320.550000 ;
      RECT 0.000000 319.750000 679.200000 320.250000 ;
      RECT 0.720000 319.450000 679.200000 319.750000 ;
      RECT 0.000000 318.950000 679.200000 319.450000 ;
      RECT 0.720000 318.650000 679.200000 318.950000 ;
      RECT 0.000000 318.150000 679.200000 318.650000 ;
      RECT 0.720000 317.850000 679.200000 318.150000 ;
      RECT 0.000000 317.350000 679.200000 317.850000 ;
      RECT 0.720000 317.050000 679.200000 317.350000 ;
      RECT 0.000000 316.550000 679.200000 317.050000 ;
      RECT 0.720000 316.250000 679.200000 316.550000 ;
      RECT 0.000000 315.750000 679.200000 316.250000 ;
      RECT 0.720000 315.450000 679.200000 315.750000 ;
      RECT 0.000000 314.950000 679.200000 315.450000 ;
      RECT 0.720000 314.650000 679.200000 314.950000 ;
      RECT 0.000000 314.150000 679.200000 314.650000 ;
      RECT 0.720000 313.850000 679.200000 314.150000 ;
      RECT 0.000000 313.350000 679.200000 313.850000 ;
      RECT 0.720000 313.050000 679.200000 313.350000 ;
      RECT 0.000000 312.550000 679.200000 313.050000 ;
      RECT 0.720000 312.250000 679.200000 312.550000 ;
      RECT 0.000000 311.750000 679.200000 312.250000 ;
      RECT 0.720000 311.450000 679.200000 311.750000 ;
      RECT 0.000000 310.950000 679.200000 311.450000 ;
      RECT 0.720000 310.650000 679.200000 310.950000 ;
      RECT 0.000000 310.150000 679.200000 310.650000 ;
      RECT 0.720000 309.850000 679.200000 310.150000 ;
      RECT 0.000000 309.350000 679.200000 309.850000 ;
      RECT 0.720000 309.050000 679.200000 309.350000 ;
      RECT 0.000000 308.550000 679.200000 309.050000 ;
      RECT 0.720000 308.250000 679.200000 308.550000 ;
      RECT 0.000000 307.750000 679.200000 308.250000 ;
      RECT 0.720000 307.450000 679.200000 307.750000 ;
      RECT 0.000000 306.950000 679.200000 307.450000 ;
      RECT 0.720000 306.650000 679.200000 306.950000 ;
      RECT 0.000000 306.150000 679.200000 306.650000 ;
      RECT 0.720000 305.850000 679.200000 306.150000 ;
      RECT 0.000000 305.350000 679.200000 305.850000 ;
      RECT 0.720000 305.050000 679.200000 305.350000 ;
      RECT 0.000000 304.550000 679.200000 305.050000 ;
      RECT 0.720000 304.250000 679.200000 304.550000 ;
      RECT 0.000000 303.750000 679.200000 304.250000 ;
      RECT 0.720000 303.450000 679.200000 303.750000 ;
      RECT 0.000000 302.950000 679.200000 303.450000 ;
      RECT 0.720000 302.650000 679.200000 302.950000 ;
      RECT 0.000000 302.150000 679.200000 302.650000 ;
      RECT 0.720000 301.850000 679.200000 302.150000 ;
      RECT 0.000000 301.350000 679.200000 301.850000 ;
      RECT 0.720000 301.050000 679.200000 301.350000 ;
      RECT 0.000000 300.550000 679.200000 301.050000 ;
      RECT 0.720000 300.250000 679.200000 300.550000 ;
      RECT 0.000000 299.750000 679.200000 300.250000 ;
      RECT 0.720000 299.450000 679.200000 299.750000 ;
      RECT 0.000000 298.950000 679.200000 299.450000 ;
      RECT 0.720000 298.650000 679.200000 298.950000 ;
      RECT 0.000000 298.150000 679.200000 298.650000 ;
      RECT 0.720000 297.850000 679.200000 298.150000 ;
      RECT 0.000000 297.350000 679.200000 297.850000 ;
      RECT 0.720000 297.050000 679.200000 297.350000 ;
      RECT 0.000000 296.550000 679.200000 297.050000 ;
      RECT 0.720000 296.250000 679.200000 296.550000 ;
      RECT 0.000000 295.750000 679.200000 296.250000 ;
      RECT 0.720000 295.450000 679.200000 295.750000 ;
      RECT 0.000000 294.950000 679.200000 295.450000 ;
      RECT 0.720000 294.650000 679.200000 294.950000 ;
      RECT 0.000000 294.150000 679.200000 294.650000 ;
      RECT 0.720000 293.850000 679.200000 294.150000 ;
      RECT 0.000000 293.350000 679.200000 293.850000 ;
      RECT 0.720000 293.050000 679.200000 293.350000 ;
      RECT 0.000000 292.550000 679.200000 293.050000 ;
      RECT 0.720000 292.250000 679.200000 292.550000 ;
      RECT 0.000000 291.750000 679.200000 292.250000 ;
      RECT 0.720000 291.450000 679.200000 291.750000 ;
      RECT 0.000000 290.950000 679.200000 291.450000 ;
      RECT 0.720000 290.650000 679.200000 290.950000 ;
      RECT 0.000000 290.150000 679.200000 290.650000 ;
      RECT 0.720000 289.850000 679.200000 290.150000 ;
      RECT 0.000000 289.350000 679.200000 289.850000 ;
      RECT 0.720000 289.050000 679.200000 289.350000 ;
      RECT 0.000000 288.550000 679.200000 289.050000 ;
      RECT 0.720000 288.250000 679.200000 288.550000 ;
      RECT 0.000000 287.750000 679.200000 288.250000 ;
      RECT 0.720000 287.450000 679.200000 287.750000 ;
      RECT 0.000000 286.950000 679.200000 287.450000 ;
      RECT 0.720000 286.650000 679.200000 286.950000 ;
      RECT 0.000000 286.150000 679.200000 286.650000 ;
      RECT 0.720000 285.850000 679.200000 286.150000 ;
      RECT 0.000000 285.350000 679.200000 285.850000 ;
      RECT 0.720000 285.050000 679.200000 285.350000 ;
      RECT 0.000000 284.550000 679.200000 285.050000 ;
      RECT 0.720000 284.250000 679.200000 284.550000 ;
      RECT 0.000000 283.750000 679.200000 284.250000 ;
      RECT 0.720000 283.450000 679.200000 283.750000 ;
      RECT 0.000000 282.950000 679.200000 283.450000 ;
      RECT 0.720000 282.650000 679.200000 282.950000 ;
      RECT 0.000000 282.150000 679.200000 282.650000 ;
      RECT 0.720000 281.850000 679.200000 282.150000 ;
      RECT 0.000000 281.350000 679.200000 281.850000 ;
      RECT 0.720000 281.050000 679.200000 281.350000 ;
      RECT 0.000000 280.550000 679.200000 281.050000 ;
      RECT 0.720000 280.250000 679.200000 280.550000 ;
      RECT 0.000000 279.750000 679.200000 280.250000 ;
      RECT 0.720000 279.450000 679.200000 279.750000 ;
      RECT 0.000000 278.950000 679.200000 279.450000 ;
      RECT 0.720000 278.650000 679.200000 278.950000 ;
      RECT 0.000000 278.150000 679.200000 278.650000 ;
      RECT 0.720000 277.850000 679.200000 278.150000 ;
      RECT 0.000000 277.350000 679.200000 277.850000 ;
      RECT 0.720000 277.050000 679.200000 277.350000 ;
      RECT 0.000000 276.550000 679.200000 277.050000 ;
      RECT 0.720000 276.250000 679.200000 276.550000 ;
      RECT 0.000000 275.750000 679.200000 276.250000 ;
      RECT 0.720000 275.450000 679.200000 275.750000 ;
      RECT 0.000000 274.950000 679.200000 275.450000 ;
      RECT 0.720000 274.650000 679.200000 274.950000 ;
      RECT 0.000000 274.150000 679.200000 274.650000 ;
      RECT 0.720000 273.850000 679.200000 274.150000 ;
      RECT 0.000000 273.350000 679.200000 273.850000 ;
      RECT 0.720000 273.050000 679.200000 273.350000 ;
      RECT 0.000000 272.550000 679.200000 273.050000 ;
      RECT 0.720000 272.250000 679.200000 272.550000 ;
      RECT 0.000000 271.750000 679.200000 272.250000 ;
      RECT 0.720000 271.450000 679.200000 271.750000 ;
      RECT 0.000000 270.950000 679.200000 271.450000 ;
      RECT 0.720000 270.650000 679.200000 270.950000 ;
      RECT 0.000000 270.150000 679.200000 270.650000 ;
      RECT 0.720000 269.850000 679.200000 270.150000 ;
      RECT 0.000000 269.350000 679.200000 269.850000 ;
      RECT 0.720000 269.050000 679.200000 269.350000 ;
      RECT 0.000000 268.550000 679.200000 269.050000 ;
      RECT 0.720000 268.250000 679.200000 268.550000 ;
      RECT 0.000000 267.750000 679.200000 268.250000 ;
      RECT 0.720000 267.450000 679.200000 267.750000 ;
      RECT 0.000000 266.950000 679.200000 267.450000 ;
      RECT 0.720000 266.650000 679.200000 266.950000 ;
      RECT 0.000000 266.150000 679.200000 266.650000 ;
      RECT 0.720000 265.850000 679.200000 266.150000 ;
      RECT 0.000000 265.350000 679.200000 265.850000 ;
      RECT 0.720000 265.050000 679.200000 265.350000 ;
      RECT 0.000000 264.550000 679.200000 265.050000 ;
      RECT 0.720000 264.250000 679.200000 264.550000 ;
      RECT 0.000000 263.750000 679.200000 264.250000 ;
      RECT 0.720000 263.450000 679.200000 263.750000 ;
      RECT 0.000000 0.760000 679.200000 263.450000 ;
      RECT 390.510000 0.000000 679.200000 0.760000 ;
      RECT 389.710000 0.000000 390.090000 0.760000 ;
      RECT 388.910000 0.000000 389.290000 0.760000 ;
      RECT 388.110000 0.000000 388.490000 0.760000 ;
      RECT 387.310000 0.000000 387.690000 0.760000 ;
      RECT 386.510000 0.000000 386.890000 0.760000 ;
      RECT 385.710000 0.000000 386.090000 0.760000 ;
      RECT 384.910000 0.000000 385.290000 0.760000 ;
      RECT 384.110000 0.000000 384.490000 0.760000 ;
      RECT 383.310000 0.000000 383.690000 0.760000 ;
      RECT 382.510000 0.000000 382.890000 0.760000 ;
      RECT 381.710000 0.000000 382.090000 0.760000 ;
      RECT 380.910000 0.000000 381.290000 0.760000 ;
      RECT 380.110000 0.000000 380.490000 0.760000 ;
      RECT 379.310000 0.000000 379.690000 0.760000 ;
      RECT 378.510000 0.000000 378.890000 0.760000 ;
      RECT 377.710000 0.000000 378.090000 0.760000 ;
      RECT 376.910000 0.000000 377.290000 0.760000 ;
      RECT 376.110000 0.000000 376.490000 0.760000 ;
      RECT 375.310000 0.000000 375.690000 0.760000 ;
      RECT 374.510000 0.000000 374.890000 0.760000 ;
      RECT 373.710000 0.000000 374.090000 0.760000 ;
      RECT 372.910000 0.000000 373.290000 0.760000 ;
      RECT 372.110000 0.000000 372.490000 0.760000 ;
      RECT 371.310000 0.000000 371.690000 0.760000 ;
      RECT 370.510000 0.000000 370.890000 0.760000 ;
      RECT 369.710000 0.000000 370.090000 0.760000 ;
      RECT 368.910000 0.000000 369.290000 0.760000 ;
      RECT 368.110000 0.000000 368.490000 0.760000 ;
      RECT 367.310000 0.000000 367.690000 0.760000 ;
      RECT 366.510000 0.000000 366.890000 0.760000 ;
      RECT 365.710000 0.000000 366.090000 0.760000 ;
      RECT 364.910000 0.000000 365.290000 0.760000 ;
      RECT 364.110000 0.000000 364.490000 0.760000 ;
      RECT 363.310000 0.000000 363.690000 0.760000 ;
      RECT 362.510000 0.000000 362.890000 0.760000 ;
      RECT 361.710000 0.000000 362.090000 0.760000 ;
      RECT 360.910000 0.000000 361.290000 0.760000 ;
      RECT 360.110000 0.000000 360.490000 0.760000 ;
      RECT 359.310000 0.000000 359.690000 0.760000 ;
      RECT 358.510000 0.000000 358.890000 0.760000 ;
      RECT 357.710000 0.000000 358.090000 0.760000 ;
      RECT 356.910000 0.000000 357.290000 0.760000 ;
      RECT 356.110000 0.000000 356.490000 0.760000 ;
      RECT 355.310000 0.000000 355.690000 0.760000 ;
      RECT 354.510000 0.000000 354.890000 0.760000 ;
      RECT 353.710000 0.000000 354.090000 0.760000 ;
      RECT 352.910000 0.000000 353.290000 0.760000 ;
      RECT 352.110000 0.000000 352.490000 0.760000 ;
      RECT 351.310000 0.000000 351.690000 0.760000 ;
      RECT 350.510000 0.000000 350.890000 0.760000 ;
      RECT 349.710000 0.000000 350.090000 0.760000 ;
      RECT 348.910000 0.000000 349.290000 0.760000 ;
      RECT 348.110000 0.000000 348.490000 0.760000 ;
      RECT 347.310000 0.000000 347.690000 0.760000 ;
      RECT 346.510000 0.000000 346.890000 0.760000 ;
      RECT 345.710000 0.000000 346.090000 0.760000 ;
      RECT 344.910000 0.000000 345.290000 0.760000 ;
      RECT 344.110000 0.000000 344.490000 0.760000 ;
      RECT 343.310000 0.000000 343.690000 0.760000 ;
      RECT 342.510000 0.000000 342.890000 0.760000 ;
      RECT 341.710000 0.000000 342.090000 0.760000 ;
      RECT 340.910000 0.000000 341.290000 0.760000 ;
      RECT 340.110000 0.000000 340.490000 0.760000 ;
      RECT 339.310000 0.000000 339.690000 0.760000 ;
      RECT 338.510000 0.000000 338.890000 0.760000 ;
      RECT 337.710000 0.000000 338.090000 0.760000 ;
      RECT 336.910000 0.000000 337.290000 0.760000 ;
      RECT 336.110000 0.000000 336.490000 0.760000 ;
      RECT 335.310000 0.000000 335.690000 0.760000 ;
      RECT 334.510000 0.000000 334.890000 0.760000 ;
      RECT 333.710000 0.000000 334.090000 0.760000 ;
      RECT 332.910000 0.000000 333.290000 0.760000 ;
      RECT 332.110000 0.000000 332.490000 0.760000 ;
      RECT 331.310000 0.000000 331.690000 0.760000 ;
      RECT 330.510000 0.000000 330.890000 0.760000 ;
      RECT 329.710000 0.000000 330.090000 0.760000 ;
      RECT 328.910000 0.000000 329.290000 0.760000 ;
      RECT 328.110000 0.000000 328.490000 0.760000 ;
      RECT 327.310000 0.000000 327.690000 0.760000 ;
      RECT 326.510000 0.000000 326.890000 0.760000 ;
      RECT 325.710000 0.000000 326.090000 0.760000 ;
      RECT 324.910000 0.000000 325.290000 0.760000 ;
      RECT 324.110000 0.000000 324.490000 0.760000 ;
      RECT 323.310000 0.000000 323.690000 0.760000 ;
      RECT 322.510000 0.000000 322.890000 0.760000 ;
      RECT 321.710000 0.000000 322.090000 0.760000 ;
      RECT 320.910000 0.000000 321.290000 0.760000 ;
      RECT 320.110000 0.000000 320.490000 0.760000 ;
      RECT 319.310000 0.000000 319.690000 0.760000 ;
      RECT 318.510000 0.000000 318.890000 0.760000 ;
      RECT 317.710000 0.000000 318.090000 0.760000 ;
      RECT 316.910000 0.000000 317.290000 0.760000 ;
      RECT 316.110000 0.000000 316.490000 0.760000 ;
      RECT 315.310000 0.000000 315.690000 0.760000 ;
      RECT 314.510000 0.000000 314.890000 0.760000 ;
      RECT 313.710000 0.000000 314.090000 0.760000 ;
      RECT 312.910000 0.000000 313.290000 0.760000 ;
      RECT 312.110000 0.000000 312.490000 0.760000 ;
      RECT 311.310000 0.000000 311.690000 0.760000 ;
      RECT 310.510000 0.000000 310.890000 0.760000 ;
      RECT 309.710000 0.000000 310.090000 0.760000 ;
      RECT 308.910000 0.000000 309.290000 0.760000 ;
      RECT 308.110000 0.000000 308.490000 0.760000 ;
      RECT 307.310000 0.000000 307.690000 0.760000 ;
      RECT 306.510000 0.000000 306.890000 0.760000 ;
      RECT 305.710000 0.000000 306.090000 0.760000 ;
      RECT 304.910000 0.000000 305.290000 0.760000 ;
      RECT 304.110000 0.000000 304.490000 0.760000 ;
      RECT 303.310000 0.000000 303.690000 0.760000 ;
      RECT 302.510000 0.000000 302.890000 0.760000 ;
      RECT 301.710000 0.000000 302.090000 0.760000 ;
      RECT 300.910000 0.000000 301.290000 0.760000 ;
      RECT 300.110000 0.000000 300.490000 0.760000 ;
      RECT 299.310000 0.000000 299.690000 0.760000 ;
      RECT 298.510000 0.000000 298.890000 0.760000 ;
      RECT 297.710000 0.000000 298.090000 0.760000 ;
      RECT 296.910000 0.000000 297.290000 0.760000 ;
      RECT 296.110000 0.000000 296.490000 0.760000 ;
      RECT 295.310000 0.000000 295.690000 0.760000 ;
      RECT 294.510000 0.000000 294.890000 0.760000 ;
      RECT 293.710000 0.000000 294.090000 0.760000 ;
      RECT 292.910000 0.000000 293.290000 0.760000 ;
      RECT 292.110000 0.000000 292.490000 0.760000 ;
      RECT 291.310000 0.000000 291.690000 0.760000 ;
      RECT 290.510000 0.000000 290.890000 0.760000 ;
      RECT 289.710000 0.000000 290.090000 0.760000 ;
      RECT 288.910000 0.000000 289.290000 0.760000 ;
      RECT 0.000000 0.000000 288.490000 0.760000 ;
    LAYER M4 ;
      RECT 0.000000 0.000000 679.200000 677.000000 ;
    LAYER M5 ;
      RECT 0.000000 0.000000 679.200000 677.000000 ;
    LAYER M6 ;
      RECT 0.000000 0.000000 679.200000 677.000000 ;
    LAYER M7 ;
      RECT 0.000000 0.000000 679.200000 677.000000 ;
    LAYER M8 ;
      RECT 0.000000 0.000000 679.200000 677.000000 ;
  END
END fullchip

END LIBRARY
