##
## LEF for PtnCells ;
## created by Innovus v19.17-s077_1 on Mon Feb 27 21:10:15 2023
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO fullchip
  CLASS BLOCK ;
  SIZE 697.600000 BY 695.000000 ;
  FOREIGN fullchip 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 288.950000 0.600000 289.050000 ;
    END
  END clk
  PIN mem_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 404.950000 0.600000 405.050000 ;
    END
  END mem_in[127]
  PIN mem_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 404.150000 0.600000 404.250000 ;
    END
  END mem_in[126]
  PIN mem_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 403.350000 0.600000 403.450000 ;
    END
  END mem_in[125]
  PIN mem_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 402.550000 0.600000 402.650000 ;
    END
  END mem_in[124]
  PIN mem_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 401.750000 0.600000 401.850000 ;
    END
  END mem_in[123]
  PIN mem_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 400.950000 0.600000 401.050000 ;
    END
  END mem_in[122]
  PIN mem_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 400.150000 0.600000 400.250000 ;
    END
  END mem_in[121]
  PIN mem_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 399.350000 0.600000 399.450000 ;
    END
  END mem_in[120]
  PIN mem_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 398.550000 0.600000 398.650000 ;
    END
  END mem_in[119]
  PIN mem_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 397.750000 0.600000 397.850000 ;
    END
  END mem_in[118]
  PIN mem_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 396.950000 0.600000 397.050000 ;
    END
  END mem_in[117]
  PIN mem_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 396.150000 0.600000 396.250000 ;
    END
  END mem_in[116]
  PIN mem_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 395.350000 0.600000 395.450000 ;
    END
  END mem_in[115]
  PIN mem_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 394.550000 0.600000 394.650000 ;
    END
  END mem_in[114]
  PIN mem_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 393.750000 0.600000 393.850000 ;
    END
  END mem_in[113]
  PIN mem_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 392.950000 0.600000 393.050000 ;
    END
  END mem_in[112]
  PIN mem_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 392.150000 0.600000 392.250000 ;
    END
  END mem_in[111]
  PIN mem_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 391.350000 0.600000 391.450000 ;
    END
  END mem_in[110]
  PIN mem_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 390.550000 0.600000 390.650000 ;
    END
  END mem_in[109]
  PIN mem_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 389.750000 0.600000 389.850000 ;
    END
  END mem_in[108]
  PIN mem_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 388.950000 0.600000 389.050000 ;
    END
  END mem_in[107]
  PIN mem_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 388.150000 0.600000 388.250000 ;
    END
  END mem_in[106]
  PIN mem_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 387.350000 0.600000 387.450000 ;
    END
  END mem_in[105]
  PIN mem_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 386.550000 0.600000 386.650000 ;
    END
  END mem_in[104]
  PIN mem_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 385.750000 0.600000 385.850000 ;
    END
  END mem_in[103]
  PIN mem_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 384.950000 0.600000 385.050000 ;
    END
  END mem_in[102]
  PIN mem_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 384.150000 0.600000 384.250000 ;
    END
  END mem_in[101]
  PIN mem_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 383.350000 0.600000 383.450000 ;
    END
  END mem_in[100]
  PIN mem_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 382.550000 0.600000 382.650000 ;
    END
  END mem_in[99]
  PIN mem_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 381.750000 0.600000 381.850000 ;
    END
  END mem_in[98]
  PIN mem_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 380.950000 0.600000 381.050000 ;
    END
  END mem_in[97]
  PIN mem_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 380.150000 0.600000 380.250000 ;
    END
  END mem_in[96]
  PIN mem_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 379.350000 0.600000 379.450000 ;
    END
  END mem_in[95]
  PIN mem_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 378.550000 0.600000 378.650000 ;
    END
  END mem_in[94]
  PIN mem_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 377.750000 0.600000 377.850000 ;
    END
  END mem_in[93]
  PIN mem_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 376.950000 0.600000 377.050000 ;
    END
  END mem_in[92]
  PIN mem_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 376.150000 0.600000 376.250000 ;
    END
  END mem_in[91]
  PIN mem_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 375.350000 0.600000 375.450000 ;
    END
  END mem_in[90]
  PIN mem_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 374.550000 0.600000 374.650000 ;
    END
  END mem_in[89]
  PIN mem_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 373.750000 0.600000 373.850000 ;
    END
  END mem_in[88]
  PIN mem_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 372.950000 0.600000 373.050000 ;
    END
  END mem_in[87]
  PIN mem_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 372.150000 0.600000 372.250000 ;
    END
  END mem_in[86]
  PIN mem_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 371.350000 0.600000 371.450000 ;
    END
  END mem_in[85]
  PIN mem_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 370.550000 0.600000 370.650000 ;
    END
  END mem_in[84]
  PIN mem_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 369.750000 0.600000 369.850000 ;
    END
  END mem_in[83]
  PIN mem_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 368.950000 0.600000 369.050000 ;
    END
  END mem_in[82]
  PIN mem_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 368.150000 0.600000 368.250000 ;
    END
  END mem_in[81]
  PIN mem_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 367.350000 0.600000 367.450000 ;
    END
  END mem_in[80]
  PIN mem_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 366.550000 0.600000 366.650000 ;
    END
  END mem_in[79]
  PIN mem_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 365.750000 0.600000 365.850000 ;
    END
  END mem_in[78]
  PIN mem_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 364.950000 0.600000 365.050000 ;
    END
  END mem_in[77]
  PIN mem_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 364.150000 0.600000 364.250000 ;
    END
  END mem_in[76]
  PIN mem_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 363.350000 0.600000 363.450000 ;
    END
  END mem_in[75]
  PIN mem_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 362.550000 0.600000 362.650000 ;
    END
  END mem_in[74]
  PIN mem_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 361.750000 0.600000 361.850000 ;
    END
  END mem_in[73]
  PIN mem_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 360.950000 0.600000 361.050000 ;
    END
  END mem_in[72]
  PIN mem_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 360.150000 0.600000 360.250000 ;
    END
  END mem_in[71]
  PIN mem_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 359.350000 0.600000 359.450000 ;
    END
  END mem_in[70]
  PIN mem_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 358.550000 0.600000 358.650000 ;
    END
  END mem_in[69]
  PIN mem_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 357.750000 0.600000 357.850000 ;
    END
  END mem_in[68]
  PIN mem_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 356.950000 0.600000 357.050000 ;
    END
  END mem_in[67]
  PIN mem_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 356.150000 0.600000 356.250000 ;
    END
  END mem_in[66]
  PIN mem_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 355.350000 0.600000 355.450000 ;
    END
  END mem_in[65]
  PIN mem_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 354.550000 0.600000 354.650000 ;
    END
  END mem_in[64]
  PIN mem_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 353.750000 0.600000 353.850000 ;
    END
  END mem_in[63]
  PIN mem_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 352.950000 0.600000 353.050000 ;
    END
  END mem_in[62]
  PIN mem_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 352.150000 0.600000 352.250000 ;
    END
  END mem_in[61]
  PIN mem_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 351.350000 0.600000 351.450000 ;
    END
  END mem_in[60]
  PIN mem_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 350.550000 0.600000 350.650000 ;
    END
  END mem_in[59]
  PIN mem_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 349.750000 0.600000 349.850000 ;
    END
  END mem_in[58]
  PIN mem_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 348.950000 0.600000 349.050000 ;
    END
  END mem_in[57]
  PIN mem_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 348.150000 0.600000 348.250000 ;
    END
  END mem_in[56]
  PIN mem_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 347.350000 0.600000 347.450000 ;
    END
  END mem_in[55]
  PIN mem_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 346.550000 0.600000 346.650000 ;
    END
  END mem_in[54]
  PIN mem_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 345.750000 0.600000 345.850000 ;
    END
  END mem_in[53]
  PIN mem_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 344.950000 0.600000 345.050000 ;
    END
  END mem_in[52]
  PIN mem_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 344.150000 0.600000 344.250000 ;
    END
  END mem_in[51]
  PIN mem_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 343.350000 0.600000 343.450000 ;
    END
  END mem_in[50]
  PIN mem_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 342.550000 0.600000 342.650000 ;
    END
  END mem_in[49]
  PIN mem_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 341.750000 0.600000 341.850000 ;
    END
  END mem_in[48]
  PIN mem_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 340.950000 0.600000 341.050000 ;
    END
  END mem_in[47]
  PIN mem_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 340.150000 0.600000 340.250000 ;
    END
  END mem_in[46]
  PIN mem_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 339.350000 0.600000 339.450000 ;
    END
  END mem_in[45]
  PIN mem_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 338.550000 0.600000 338.650000 ;
    END
  END mem_in[44]
  PIN mem_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 337.750000 0.600000 337.850000 ;
    END
  END mem_in[43]
  PIN mem_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 336.950000 0.600000 337.050000 ;
    END
  END mem_in[42]
  PIN mem_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 336.150000 0.600000 336.250000 ;
    END
  END mem_in[41]
  PIN mem_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 335.350000 0.600000 335.450000 ;
    END
  END mem_in[40]
  PIN mem_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 334.550000 0.600000 334.650000 ;
    END
  END mem_in[39]
  PIN mem_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 333.750000 0.600000 333.850000 ;
    END
  END mem_in[38]
  PIN mem_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 332.950000 0.600000 333.050000 ;
    END
  END mem_in[37]
  PIN mem_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 332.150000 0.600000 332.250000 ;
    END
  END mem_in[36]
  PIN mem_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 331.350000 0.600000 331.450000 ;
    END
  END mem_in[35]
  PIN mem_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 330.550000 0.600000 330.650000 ;
    END
  END mem_in[34]
  PIN mem_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 329.750000 0.600000 329.850000 ;
    END
  END mem_in[33]
  PIN mem_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 328.950000 0.600000 329.050000 ;
    END
  END mem_in[32]
  PIN mem_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 328.150000 0.600000 328.250000 ;
    END
  END mem_in[31]
  PIN mem_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 327.350000 0.600000 327.450000 ;
    END
  END mem_in[30]
  PIN mem_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 326.550000 0.600000 326.650000 ;
    END
  END mem_in[29]
  PIN mem_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 325.750000 0.600000 325.850000 ;
    END
  END mem_in[28]
  PIN mem_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 324.950000 0.600000 325.050000 ;
    END
  END mem_in[27]
  PIN mem_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 324.150000 0.600000 324.250000 ;
    END
  END mem_in[26]
  PIN mem_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 323.350000 0.600000 323.450000 ;
    END
  END mem_in[25]
  PIN mem_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 322.550000 0.600000 322.650000 ;
    END
  END mem_in[24]
  PIN mem_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 321.750000 0.600000 321.850000 ;
    END
  END mem_in[23]
  PIN mem_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 320.950000 0.600000 321.050000 ;
    END
  END mem_in[22]
  PIN mem_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 320.150000 0.600000 320.250000 ;
    END
  END mem_in[21]
  PIN mem_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 319.350000 0.600000 319.450000 ;
    END
  END mem_in[20]
  PIN mem_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 318.550000 0.600000 318.650000 ;
    END
  END mem_in[19]
  PIN mem_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 317.750000 0.600000 317.850000 ;
    END
  END mem_in[18]
  PIN mem_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 316.950000 0.600000 317.050000 ;
    END
  END mem_in[17]
  PIN mem_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 316.150000 0.600000 316.250000 ;
    END
  END mem_in[16]
  PIN mem_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 315.350000 0.600000 315.450000 ;
    END
  END mem_in[15]
  PIN mem_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 314.550000 0.600000 314.650000 ;
    END
  END mem_in[14]
  PIN mem_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 313.750000 0.600000 313.850000 ;
    END
  END mem_in[13]
  PIN mem_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 312.950000 0.600000 313.050000 ;
    END
  END mem_in[12]
  PIN mem_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 312.150000 0.600000 312.250000 ;
    END
  END mem_in[11]
  PIN mem_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 311.350000 0.600000 311.450000 ;
    END
  END mem_in[10]
  PIN mem_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 310.550000 0.600000 310.650000 ;
    END
  END mem_in[9]
  PIN mem_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 309.750000 0.600000 309.850000 ;
    END
  END mem_in[8]
  PIN mem_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 308.950000 0.600000 309.050000 ;
    END
  END mem_in[7]
  PIN mem_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 308.150000 0.600000 308.250000 ;
    END
  END mem_in[6]
  PIN mem_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 307.350000 0.600000 307.450000 ;
    END
  END mem_in[5]
  PIN mem_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 306.550000 0.600000 306.650000 ;
    END
  END mem_in[4]
  PIN mem_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 305.750000 0.600000 305.850000 ;
    END
  END mem_in[3]
  PIN mem_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 304.950000 0.600000 305.050000 ;
    END
  END mem_in[2]
  PIN mem_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 304.150000 0.600000 304.250000 ;
    END
  END mem_in[1]
  PIN mem_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 303.350000 0.600000 303.450000 ;
    END
  END mem_in[0]
  PIN inst[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 302.550000 0.600000 302.650000 ;
    END
  END inst[16]
  PIN inst[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 301.750000 0.600000 301.850000 ;
    END
  END inst[15]
  PIN inst[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 300.950000 0.600000 301.050000 ;
    END
  END inst[14]
  PIN inst[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 300.150000 0.600000 300.250000 ;
    END
  END inst[13]
  PIN inst[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 299.350000 0.600000 299.450000 ;
    END
  END inst[12]
  PIN inst[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 298.550000 0.600000 298.650000 ;
    END
  END inst[11]
  PIN inst[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 297.750000 0.600000 297.850000 ;
    END
  END inst[10]
  PIN inst[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 296.950000 0.600000 297.050000 ;
    END
  END inst[9]
  PIN inst[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 296.150000 0.600000 296.250000 ;
    END
  END inst[8]
  PIN inst[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 295.350000 0.600000 295.450000 ;
    END
  END inst[7]
  PIN inst[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 294.550000 0.600000 294.650000 ;
    END
  END inst[6]
  PIN inst[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 293.750000 0.600000 293.850000 ;
    END
  END inst[5]
  PIN inst[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 292.950000 0.600000 293.050000 ;
    END
  END inst[4]
  PIN inst[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 292.150000 0.600000 292.250000 ;
    END
  END inst[3]
  PIN inst[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 291.350000 0.600000 291.450000 ;
    END
  END inst[2]
  PIN inst[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 290.550000 0.600000 290.650000 ;
    END
  END inst[1]
  PIN inst[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 289.750000 0.600000 289.850000 ;
    END
  END inst[0]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 405.750000 0.600000 405.850000 ;
    END
  END reset
  PIN sum_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 275.650000 0.000000 275.750000 0.600000 ;
    END
  END sum_out[23]
  PIN sum_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 276.450000 0.000000 276.550000 0.600000 ;
    END
  END sum_out[22]
  PIN sum_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 277.250000 0.000000 277.350000 0.600000 ;
    END
  END sum_out[21]
  PIN sum_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 278.050000 0.000000 278.150000 0.600000 ;
    END
  END sum_out[20]
  PIN sum_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 278.850000 0.000000 278.950000 0.600000 ;
    END
  END sum_out[19]
  PIN sum_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 279.650000 0.000000 279.750000 0.600000 ;
    END
  END sum_out[18]
  PIN sum_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 280.450000 0.000000 280.550000 0.600000 ;
    END
  END sum_out[17]
  PIN sum_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 281.250000 0.000000 281.350000 0.600000 ;
    END
  END sum_out[16]
  PIN sum_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 282.050000 0.000000 282.150000 0.600000 ;
    END
  END sum_out[15]
  PIN sum_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 282.850000 0.000000 282.950000 0.600000 ;
    END
  END sum_out[14]
  PIN sum_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 283.650000 0.000000 283.750000 0.600000 ;
    END
  END sum_out[13]
  PIN sum_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 284.450000 0.000000 284.550000 0.600000 ;
    END
  END sum_out[12]
  PIN sum_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 285.250000 0.000000 285.350000 0.600000 ;
    END
  END sum_out[11]
  PIN sum_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 286.050000 0.000000 286.150000 0.600000 ;
    END
  END sum_out[10]
  PIN sum_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 286.850000 0.000000 286.950000 0.600000 ;
    END
  END sum_out[9]
  PIN sum_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 287.650000 0.000000 287.750000 0.600000 ;
    END
  END sum_out[8]
  PIN sum_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 288.450000 0.000000 288.550000 0.600000 ;
    END
  END sum_out[7]
  PIN sum_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 289.250000 0.000000 289.350000 0.600000 ;
    END
  END sum_out[6]
  PIN sum_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 290.050000 0.000000 290.150000 0.600000 ;
    END
  END sum_out[5]
  PIN sum_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 290.850000 0.000000 290.950000 0.600000 ;
    END
  END sum_out[4]
  PIN sum_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 291.650000 0.000000 291.750000 0.600000 ;
    END
  END sum_out[3]
  PIN sum_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 292.450000 0.000000 292.550000 0.600000 ;
    END
  END sum_out[2]
  PIN sum_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 293.250000 0.000000 293.350000 0.600000 ;
    END
  END sum_out[1]
  PIN sum_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 294.050000 0.000000 294.150000 0.600000 ;
    END
  END sum_out[0]
  PIN out[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 294.850000 0.000000 294.950000 0.600000 ;
    END
  END out[159]
  PIN out[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 295.650000 0.000000 295.750000 0.600000 ;
    END
  END out[158]
  PIN out[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 296.450000 0.000000 296.550000 0.600000 ;
    END
  END out[157]
  PIN out[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 297.250000 0.000000 297.350000 0.600000 ;
    END
  END out[156]
  PIN out[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 298.050000 0.000000 298.150000 0.600000 ;
    END
  END out[155]
  PIN out[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 298.850000 0.000000 298.950000 0.600000 ;
    END
  END out[154]
  PIN out[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 299.650000 0.000000 299.750000 0.600000 ;
    END
  END out[153]
  PIN out[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 300.450000 0.000000 300.550000 0.600000 ;
    END
  END out[152]
  PIN out[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 301.250000 0.000000 301.350000 0.600000 ;
    END
  END out[151]
  PIN out[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 302.050000 0.000000 302.150000 0.600000 ;
    END
  END out[150]
  PIN out[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 302.850000 0.000000 302.950000 0.600000 ;
    END
  END out[149]
  PIN out[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 303.650000 0.000000 303.750000 0.600000 ;
    END
  END out[148]
  PIN out[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 304.450000 0.000000 304.550000 0.600000 ;
    END
  END out[147]
  PIN out[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 305.250000 0.000000 305.350000 0.600000 ;
    END
  END out[146]
  PIN out[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 306.050000 0.000000 306.150000 0.600000 ;
    END
  END out[145]
  PIN out[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 306.850000 0.000000 306.950000 0.600000 ;
    END
  END out[144]
  PIN out[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 307.650000 0.000000 307.750000 0.600000 ;
    END
  END out[143]
  PIN out[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 308.450000 0.000000 308.550000 0.600000 ;
    END
  END out[142]
  PIN out[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 309.250000 0.000000 309.350000 0.600000 ;
    END
  END out[141]
  PIN out[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 310.050000 0.000000 310.150000 0.600000 ;
    END
  END out[140]
  PIN out[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 310.850000 0.000000 310.950000 0.600000 ;
    END
  END out[139]
  PIN out[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 311.650000 0.000000 311.750000 0.600000 ;
    END
  END out[138]
  PIN out[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 312.450000 0.000000 312.550000 0.600000 ;
    END
  END out[137]
  PIN out[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 313.250000 0.000000 313.350000 0.600000 ;
    END
  END out[136]
  PIN out[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 314.050000 0.000000 314.150000 0.600000 ;
    END
  END out[135]
  PIN out[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 314.850000 0.000000 314.950000 0.600000 ;
    END
  END out[134]
  PIN out[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 315.650000 0.000000 315.750000 0.600000 ;
    END
  END out[133]
  PIN out[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 316.450000 0.000000 316.550000 0.600000 ;
    END
  END out[132]
  PIN out[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 317.250000 0.000000 317.350000 0.600000 ;
    END
  END out[131]
  PIN out[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 318.050000 0.000000 318.150000 0.600000 ;
    END
  END out[130]
  PIN out[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 318.850000 0.000000 318.950000 0.600000 ;
    END
  END out[129]
  PIN out[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 319.650000 0.000000 319.750000 0.600000 ;
    END
  END out[128]
  PIN out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 320.450000 0.000000 320.550000 0.600000 ;
    END
  END out[127]
  PIN out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 321.250000 0.000000 321.350000 0.600000 ;
    END
  END out[126]
  PIN out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 322.050000 0.000000 322.150000 0.600000 ;
    END
  END out[125]
  PIN out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 322.850000 0.000000 322.950000 0.600000 ;
    END
  END out[124]
  PIN out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 323.650000 0.000000 323.750000 0.600000 ;
    END
  END out[123]
  PIN out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 324.450000 0.000000 324.550000 0.600000 ;
    END
  END out[122]
  PIN out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 325.250000 0.000000 325.350000 0.600000 ;
    END
  END out[121]
  PIN out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 326.050000 0.000000 326.150000 0.600000 ;
    END
  END out[120]
  PIN out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 326.850000 0.000000 326.950000 0.600000 ;
    END
  END out[119]
  PIN out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 327.650000 0.000000 327.750000 0.600000 ;
    END
  END out[118]
  PIN out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 328.450000 0.000000 328.550000 0.600000 ;
    END
  END out[117]
  PIN out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 329.250000 0.000000 329.350000 0.600000 ;
    END
  END out[116]
  PIN out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 330.050000 0.000000 330.150000 0.600000 ;
    END
  END out[115]
  PIN out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 330.850000 0.000000 330.950000 0.600000 ;
    END
  END out[114]
  PIN out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 331.650000 0.000000 331.750000 0.600000 ;
    END
  END out[113]
  PIN out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 332.450000 0.000000 332.550000 0.600000 ;
    END
  END out[112]
  PIN out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 333.250000 0.000000 333.350000 0.600000 ;
    END
  END out[111]
  PIN out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 334.050000 0.000000 334.150000 0.600000 ;
    END
  END out[110]
  PIN out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 334.850000 0.000000 334.950000 0.600000 ;
    END
  END out[109]
  PIN out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 335.650000 0.000000 335.750000 0.600000 ;
    END
  END out[108]
  PIN out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 336.450000 0.000000 336.550000 0.600000 ;
    END
  END out[107]
  PIN out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 337.250000 0.000000 337.350000 0.600000 ;
    END
  END out[106]
  PIN out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 338.050000 0.000000 338.150000 0.600000 ;
    END
  END out[105]
  PIN out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 338.850000 0.000000 338.950000 0.600000 ;
    END
  END out[104]
  PIN out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 339.650000 0.000000 339.750000 0.600000 ;
    END
  END out[103]
  PIN out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 340.450000 0.000000 340.550000 0.600000 ;
    END
  END out[102]
  PIN out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 341.250000 0.000000 341.350000 0.600000 ;
    END
  END out[101]
  PIN out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 342.050000 0.000000 342.150000 0.600000 ;
    END
  END out[100]
  PIN out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 342.850000 0.000000 342.950000 0.600000 ;
    END
  END out[99]
  PIN out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 343.650000 0.000000 343.750000 0.600000 ;
    END
  END out[98]
  PIN out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 344.450000 0.000000 344.550000 0.600000 ;
    END
  END out[97]
  PIN out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 345.250000 0.000000 345.350000 0.600000 ;
    END
  END out[96]
  PIN out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 346.050000 0.000000 346.150000 0.600000 ;
    END
  END out[95]
  PIN out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 346.850000 0.000000 346.950000 0.600000 ;
    END
  END out[94]
  PIN out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 347.650000 0.000000 347.750000 0.600000 ;
    END
  END out[93]
  PIN out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 348.450000 0.000000 348.550000 0.600000 ;
    END
  END out[92]
  PIN out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 349.250000 0.000000 349.350000 0.600000 ;
    END
  END out[91]
  PIN out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 350.050000 0.000000 350.150000 0.600000 ;
    END
  END out[90]
  PIN out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 350.850000 0.000000 350.950000 0.600000 ;
    END
  END out[89]
  PIN out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 351.650000 0.000000 351.750000 0.600000 ;
    END
  END out[88]
  PIN out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 352.450000 0.000000 352.550000 0.600000 ;
    END
  END out[87]
  PIN out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 353.250000 0.000000 353.350000 0.600000 ;
    END
  END out[86]
  PIN out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 354.050000 0.000000 354.150000 0.600000 ;
    END
  END out[85]
  PIN out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 354.850000 0.000000 354.950000 0.600000 ;
    END
  END out[84]
  PIN out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 355.650000 0.000000 355.750000 0.600000 ;
    END
  END out[83]
  PIN out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 356.450000 0.000000 356.550000 0.600000 ;
    END
  END out[82]
  PIN out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 357.250000 0.000000 357.350000 0.600000 ;
    END
  END out[81]
  PIN out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 358.050000 0.000000 358.150000 0.600000 ;
    END
  END out[80]
  PIN out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 358.850000 0.000000 358.950000 0.600000 ;
    END
  END out[79]
  PIN out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 359.650000 0.000000 359.750000 0.600000 ;
    END
  END out[78]
  PIN out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 360.450000 0.000000 360.550000 0.600000 ;
    END
  END out[77]
  PIN out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 361.250000 0.000000 361.350000 0.600000 ;
    END
  END out[76]
  PIN out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 362.050000 0.000000 362.150000 0.600000 ;
    END
  END out[75]
  PIN out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 362.850000 0.000000 362.950000 0.600000 ;
    END
  END out[74]
  PIN out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 363.650000 0.000000 363.750000 0.600000 ;
    END
  END out[73]
  PIN out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 364.450000 0.000000 364.550000 0.600000 ;
    END
  END out[72]
  PIN out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 365.250000 0.000000 365.350000 0.600000 ;
    END
  END out[71]
  PIN out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 366.050000 0.000000 366.150000 0.600000 ;
    END
  END out[70]
  PIN out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 366.850000 0.000000 366.950000 0.600000 ;
    END
  END out[69]
  PIN out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 367.650000 0.000000 367.750000 0.600000 ;
    END
  END out[68]
  PIN out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 368.450000 0.000000 368.550000 0.600000 ;
    END
  END out[67]
  PIN out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 369.250000 0.000000 369.350000 0.600000 ;
    END
  END out[66]
  PIN out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 370.050000 0.000000 370.150000 0.600000 ;
    END
  END out[65]
  PIN out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 370.850000 0.000000 370.950000 0.600000 ;
    END
  END out[64]
  PIN out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 371.650000 0.000000 371.750000 0.600000 ;
    END
  END out[63]
  PIN out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 372.450000 0.000000 372.550000 0.600000 ;
    END
  END out[62]
  PIN out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 373.250000 0.000000 373.350000 0.600000 ;
    END
  END out[61]
  PIN out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 374.050000 0.000000 374.150000 0.600000 ;
    END
  END out[60]
  PIN out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 374.850000 0.000000 374.950000 0.600000 ;
    END
  END out[59]
  PIN out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 375.650000 0.000000 375.750000 0.600000 ;
    END
  END out[58]
  PIN out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 376.450000 0.000000 376.550000 0.600000 ;
    END
  END out[57]
  PIN out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 377.250000 0.000000 377.350000 0.600000 ;
    END
  END out[56]
  PIN out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 378.050000 0.000000 378.150000 0.600000 ;
    END
  END out[55]
  PIN out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 378.850000 0.000000 378.950000 0.600000 ;
    END
  END out[54]
  PIN out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 379.650000 0.000000 379.750000 0.600000 ;
    END
  END out[53]
  PIN out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 380.450000 0.000000 380.550000 0.600000 ;
    END
  END out[52]
  PIN out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 381.250000 0.000000 381.350000 0.600000 ;
    END
  END out[51]
  PIN out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.050000 0.000000 382.150000 0.600000 ;
    END
  END out[50]
  PIN out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.850000 0.000000 382.950000 0.600000 ;
    END
  END out[49]
  PIN out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 383.650000 0.000000 383.750000 0.600000 ;
    END
  END out[48]
  PIN out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 384.450000 0.000000 384.550000 0.600000 ;
    END
  END out[47]
  PIN out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 385.250000 0.000000 385.350000 0.600000 ;
    END
  END out[46]
  PIN out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 386.050000 0.000000 386.150000 0.600000 ;
    END
  END out[45]
  PIN out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 386.850000 0.000000 386.950000 0.600000 ;
    END
  END out[44]
  PIN out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 387.650000 0.000000 387.750000 0.600000 ;
    END
  END out[43]
  PIN out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 388.450000 0.000000 388.550000 0.600000 ;
    END
  END out[42]
  PIN out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 389.250000 0.000000 389.350000 0.600000 ;
    END
  END out[41]
  PIN out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 390.050000 0.000000 390.150000 0.600000 ;
    END
  END out[40]
  PIN out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 390.850000 0.000000 390.950000 0.600000 ;
    END
  END out[39]
  PIN out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 391.650000 0.000000 391.750000 0.600000 ;
    END
  END out[38]
  PIN out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 392.450000 0.000000 392.550000 0.600000 ;
    END
  END out[37]
  PIN out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 393.250000 0.000000 393.350000 0.600000 ;
    END
  END out[36]
  PIN out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 394.050000 0.000000 394.150000 0.600000 ;
    END
  END out[35]
  PIN out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 394.850000 0.000000 394.950000 0.600000 ;
    END
  END out[34]
  PIN out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 395.650000 0.000000 395.750000 0.600000 ;
    END
  END out[33]
  PIN out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 396.450000 0.000000 396.550000 0.600000 ;
    END
  END out[32]
  PIN out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 397.250000 0.000000 397.350000 0.600000 ;
    END
  END out[31]
  PIN out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 398.050000 0.000000 398.150000 0.600000 ;
    END
  END out[30]
  PIN out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 398.850000 0.000000 398.950000 0.600000 ;
    END
  END out[29]
  PIN out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 399.650000 0.000000 399.750000 0.600000 ;
    END
  END out[28]
  PIN out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 400.450000 0.000000 400.550000 0.600000 ;
    END
  END out[27]
  PIN out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.250000 0.000000 401.350000 0.600000 ;
    END
  END out[26]
  PIN out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 402.050000 0.000000 402.150000 0.600000 ;
    END
  END out[25]
  PIN out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 402.850000 0.000000 402.950000 0.600000 ;
    END
  END out[24]
  PIN out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 403.650000 0.000000 403.750000 0.600000 ;
    END
  END out[23]
  PIN out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 404.450000 0.000000 404.550000 0.600000 ;
    END
  END out[22]
  PIN out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 405.250000 0.000000 405.350000 0.600000 ;
    END
  END out[21]
  PIN out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 406.050000 0.000000 406.150000 0.600000 ;
    END
  END out[20]
  PIN out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 406.850000 0.000000 406.950000 0.600000 ;
    END
  END out[19]
  PIN out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 407.650000 0.000000 407.750000 0.600000 ;
    END
  END out[18]
  PIN out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 408.450000 0.000000 408.550000 0.600000 ;
    END
  END out[17]
  PIN out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 409.250000 0.000000 409.350000 0.600000 ;
    END
  END out[16]
  PIN out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 410.050000 0.000000 410.150000 0.600000 ;
    END
  END out[15]
  PIN out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 410.850000 0.000000 410.950000 0.600000 ;
    END
  END out[14]
  PIN out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 411.650000 0.000000 411.750000 0.600000 ;
    END
  END out[13]
  PIN out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 412.450000 0.000000 412.550000 0.600000 ;
    END
  END out[12]
  PIN out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 413.250000 0.000000 413.350000 0.600000 ;
    END
  END out[11]
  PIN out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 414.050000 0.000000 414.150000 0.600000 ;
    END
  END out[10]
  PIN out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 414.850000 0.000000 414.950000 0.600000 ;
    END
  END out[9]
  PIN out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 415.650000 0.000000 415.750000 0.600000 ;
    END
  END out[8]
  PIN out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 416.450000 0.000000 416.550000 0.600000 ;
    END
  END out[7]
  PIN out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 417.250000 0.000000 417.350000 0.600000 ;
    END
  END out[6]
  PIN out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 418.050000 0.000000 418.150000 0.600000 ;
    END
  END out[5]
  PIN out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 418.850000 0.000000 418.950000 0.600000 ;
    END
  END out[4]
  PIN out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 419.650000 0.000000 419.750000 0.600000 ;
    END
  END out[3]
  PIN out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 420.450000 0.000000 420.550000 0.600000 ;
    END
  END out[2]
  PIN out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 421.250000 0.000000 421.350000 0.600000 ;
    END
  END out[1]
  PIN out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 422.050000 0.000000 422.150000 0.600000 ;
    END
  END out[0]
  OBS
    LAYER M1 ;
      RECT 0.000000 0.000000 697.600000 695.000000 ;
    LAYER M2 ;
      RECT 0.000000 0.000000 697.600000 695.000000 ;
    LAYER M3 ;
      RECT 0.000000 405.950000 697.600000 695.000000 ;
      RECT 0.720000 405.650000 697.600000 405.950000 ;
      RECT 0.000000 405.150000 697.600000 405.650000 ;
      RECT 0.720000 404.850000 697.600000 405.150000 ;
      RECT 0.000000 404.350000 697.600000 404.850000 ;
      RECT 0.720000 404.050000 697.600000 404.350000 ;
      RECT 0.000000 403.550000 697.600000 404.050000 ;
      RECT 0.720000 403.250000 697.600000 403.550000 ;
      RECT 0.000000 402.750000 697.600000 403.250000 ;
      RECT 0.720000 402.450000 697.600000 402.750000 ;
      RECT 0.000000 401.950000 697.600000 402.450000 ;
      RECT 0.720000 401.650000 697.600000 401.950000 ;
      RECT 0.000000 401.150000 697.600000 401.650000 ;
      RECT 0.720000 400.850000 697.600000 401.150000 ;
      RECT 0.000000 400.350000 697.600000 400.850000 ;
      RECT 0.720000 400.050000 697.600000 400.350000 ;
      RECT 0.000000 399.550000 697.600000 400.050000 ;
      RECT 0.720000 399.250000 697.600000 399.550000 ;
      RECT 0.000000 398.750000 697.600000 399.250000 ;
      RECT 0.720000 398.450000 697.600000 398.750000 ;
      RECT 0.000000 397.950000 697.600000 398.450000 ;
      RECT 0.720000 397.650000 697.600000 397.950000 ;
      RECT 0.000000 397.150000 697.600000 397.650000 ;
      RECT 0.720000 396.850000 697.600000 397.150000 ;
      RECT 0.000000 396.350000 697.600000 396.850000 ;
      RECT 0.720000 396.050000 697.600000 396.350000 ;
      RECT 0.000000 395.550000 697.600000 396.050000 ;
      RECT 0.720000 395.250000 697.600000 395.550000 ;
      RECT 0.000000 394.750000 697.600000 395.250000 ;
      RECT 0.720000 394.450000 697.600000 394.750000 ;
      RECT 0.000000 393.950000 697.600000 394.450000 ;
      RECT 0.720000 393.650000 697.600000 393.950000 ;
      RECT 0.000000 393.150000 697.600000 393.650000 ;
      RECT 0.720000 392.850000 697.600000 393.150000 ;
      RECT 0.000000 392.350000 697.600000 392.850000 ;
      RECT 0.720000 392.050000 697.600000 392.350000 ;
      RECT 0.000000 391.550000 697.600000 392.050000 ;
      RECT 0.720000 391.250000 697.600000 391.550000 ;
      RECT 0.000000 390.750000 697.600000 391.250000 ;
      RECT 0.720000 390.450000 697.600000 390.750000 ;
      RECT 0.000000 389.950000 697.600000 390.450000 ;
      RECT 0.720000 389.650000 697.600000 389.950000 ;
      RECT 0.000000 389.150000 697.600000 389.650000 ;
      RECT 0.720000 388.850000 697.600000 389.150000 ;
      RECT 0.000000 388.350000 697.600000 388.850000 ;
      RECT 0.720000 388.050000 697.600000 388.350000 ;
      RECT 0.000000 387.550000 697.600000 388.050000 ;
      RECT 0.720000 387.250000 697.600000 387.550000 ;
      RECT 0.000000 386.750000 697.600000 387.250000 ;
      RECT 0.720000 386.450000 697.600000 386.750000 ;
      RECT 0.000000 385.950000 697.600000 386.450000 ;
      RECT 0.720000 385.650000 697.600000 385.950000 ;
      RECT 0.000000 385.150000 697.600000 385.650000 ;
      RECT 0.720000 384.850000 697.600000 385.150000 ;
      RECT 0.000000 384.350000 697.600000 384.850000 ;
      RECT 0.720000 384.050000 697.600000 384.350000 ;
      RECT 0.000000 383.550000 697.600000 384.050000 ;
      RECT 0.720000 383.250000 697.600000 383.550000 ;
      RECT 0.000000 382.750000 697.600000 383.250000 ;
      RECT 0.720000 382.450000 697.600000 382.750000 ;
      RECT 0.000000 381.950000 697.600000 382.450000 ;
      RECT 0.720000 381.650000 697.600000 381.950000 ;
      RECT 0.000000 381.150000 697.600000 381.650000 ;
      RECT 0.720000 380.850000 697.600000 381.150000 ;
      RECT 0.000000 380.350000 697.600000 380.850000 ;
      RECT 0.720000 380.050000 697.600000 380.350000 ;
      RECT 0.000000 379.550000 697.600000 380.050000 ;
      RECT 0.720000 379.250000 697.600000 379.550000 ;
      RECT 0.000000 378.750000 697.600000 379.250000 ;
      RECT 0.720000 378.450000 697.600000 378.750000 ;
      RECT 0.000000 377.950000 697.600000 378.450000 ;
      RECT 0.720000 377.650000 697.600000 377.950000 ;
      RECT 0.000000 377.150000 697.600000 377.650000 ;
      RECT 0.720000 376.850000 697.600000 377.150000 ;
      RECT 0.000000 376.350000 697.600000 376.850000 ;
      RECT 0.720000 376.050000 697.600000 376.350000 ;
      RECT 0.000000 375.550000 697.600000 376.050000 ;
      RECT 0.720000 375.250000 697.600000 375.550000 ;
      RECT 0.000000 374.750000 697.600000 375.250000 ;
      RECT 0.720000 374.450000 697.600000 374.750000 ;
      RECT 0.000000 373.950000 697.600000 374.450000 ;
      RECT 0.720000 373.650000 697.600000 373.950000 ;
      RECT 0.000000 373.150000 697.600000 373.650000 ;
      RECT 0.720000 372.850000 697.600000 373.150000 ;
      RECT 0.000000 372.350000 697.600000 372.850000 ;
      RECT 0.720000 372.050000 697.600000 372.350000 ;
      RECT 0.000000 371.550000 697.600000 372.050000 ;
      RECT 0.720000 371.250000 697.600000 371.550000 ;
      RECT 0.000000 370.750000 697.600000 371.250000 ;
      RECT 0.720000 370.450000 697.600000 370.750000 ;
      RECT 0.000000 369.950000 697.600000 370.450000 ;
      RECT 0.720000 369.650000 697.600000 369.950000 ;
      RECT 0.000000 369.150000 697.600000 369.650000 ;
      RECT 0.720000 368.850000 697.600000 369.150000 ;
      RECT 0.000000 368.350000 697.600000 368.850000 ;
      RECT 0.720000 368.050000 697.600000 368.350000 ;
      RECT 0.000000 367.550000 697.600000 368.050000 ;
      RECT 0.720000 367.250000 697.600000 367.550000 ;
      RECT 0.000000 366.750000 697.600000 367.250000 ;
      RECT 0.720000 366.450000 697.600000 366.750000 ;
      RECT 0.000000 365.950000 697.600000 366.450000 ;
      RECT 0.720000 365.650000 697.600000 365.950000 ;
      RECT 0.000000 365.150000 697.600000 365.650000 ;
      RECT 0.720000 364.850000 697.600000 365.150000 ;
      RECT 0.000000 364.350000 697.600000 364.850000 ;
      RECT 0.720000 364.050000 697.600000 364.350000 ;
      RECT 0.000000 363.550000 697.600000 364.050000 ;
      RECT 0.720000 363.250000 697.600000 363.550000 ;
      RECT 0.000000 362.750000 697.600000 363.250000 ;
      RECT 0.720000 362.450000 697.600000 362.750000 ;
      RECT 0.000000 361.950000 697.600000 362.450000 ;
      RECT 0.720000 361.650000 697.600000 361.950000 ;
      RECT 0.000000 361.150000 697.600000 361.650000 ;
      RECT 0.720000 360.850000 697.600000 361.150000 ;
      RECT 0.000000 360.350000 697.600000 360.850000 ;
      RECT 0.720000 360.050000 697.600000 360.350000 ;
      RECT 0.000000 359.550000 697.600000 360.050000 ;
      RECT 0.720000 359.250000 697.600000 359.550000 ;
      RECT 0.000000 358.750000 697.600000 359.250000 ;
      RECT 0.720000 358.450000 697.600000 358.750000 ;
      RECT 0.000000 357.950000 697.600000 358.450000 ;
      RECT 0.720000 357.650000 697.600000 357.950000 ;
      RECT 0.000000 357.150000 697.600000 357.650000 ;
      RECT 0.720000 356.850000 697.600000 357.150000 ;
      RECT 0.000000 356.350000 697.600000 356.850000 ;
      RECT 0.720000 356.050000 697.600000 356.350000 ;
      RECT 0.000000 355.550000 697.600000 356.050000 ;
      RECT 0.720000 355.250000 697.600000 355.550000 ;
      RECT 0.000000 354.750000 697.600000 355.250000 ;
      RECT 0.720000 354.450000 697.600000 354.750000 ;
      RECT 0.000000 353.950000 697.600000 354.450000 ;
      RECT 0.720000 353.650000 697.600000 353.950000 ;
      RECT 0.000000 353.150000 697.600000 353.650000 ;
      RECT 0.720000 352.850000 697.600000 353.150000 ;
      RECT 0.000000 352.350000 697.600000 352.850000 ;
      RECT 0.720000 352.050000 697.600000 352.350000 ;
      RECT 0.000000 351.550000 697.600000 352.050000 ;
      RECT 0.720000 351.250000 697.600000 351.550000 ;
      RECT 0.000000 350.750000 697.600000 351.250000 ;
      RECT 0.720000 350.450000 697.600000 350.750000 ;
      RECT 0.000000 349.950000 697.600000 350.450000 ;
      RECT 0.720000 349.650000 697.600000 349.950000 ;
      RECT 0.000000 349.150000 697.600000 349.650000 ;
      RECT 0.720000 348.850000 697.600000 349.150000 ;
      RECT 0.000000 348.350000 697.600000 348.850000 ;
      RECT 0.720000 348.050000 697.600000 348.350000 ;
      RECT 0.000000 347.550000 697.600000 348.050000 ;
      RECT 0.720000 347.250000 697.600000 347.550000 ;
      RECT 0.000000 346.750000 697.600000 347.250000 ;
      RECT 0.720000 346.450000 697.600000 346.750000 ;
      RECT 0.000000 345.950000 697.600000 346.450000 ;
      RECT 0.720000 345.650000 697.600000 345.950000 ;
      RECT 0.000000 345.150000 697.600000 345.650000 ;
      RECT 0.720000 344.850000 697.600000 345.150000 ;
      RECT 0.000000 344.350000 697.600000 344.850000 ;
      RECT 0.720000 344.050000 697.600000 344.350000 ;
      RECT 0.000000 343.550000 697.600000 344.050000 ;
      RECT 0.720000 343.250000 697.600000 343.550000 ;
      RECT 0.000000 342.750000 697.600000 343.250000 ;
      RECT 0.720000 342.450000 697.600000 342.750000 ;
      RECT 0.000000 341.950000 697.600000 342.450000 ;
      RECT 0.720000 341.650000 697.600000 341.950000 ;
      RECT 0.000000 341.150000 697.600000 341.650000 ;
      RECT 0.720000 340.850000 697.600000 341.150000 ;
      RECT 0.000000 340.350000 697.600000 340.850000 ;
      RECT 0.720000 340.050000 697.600000 340.350000 ;
      RECT 0.000000 339.550000 697.600000 340.050000 ;
      RECT 0.720000 339.250000 697.600000 339.550000 ;
      RECT 0.000000 338.750000 697.600000 339.250000 ;
      RECT 0.720000 338.450000 697.600000 338.750000 ;
      RECT 0.000000 337.950000 697.600000 338.450000 ;
      RECT 0.720000 337.650000 697.600000 337.950000 ;
      RECT 0.000000 337.150000 697.600000 337.650000 ;
      RECT 0.720000 336.850000 697.600000 337.150000 ;
      RECT 0.000000 336.350000 697.600000 336.850000 ;
      RECT 0.720000 336.050000 697.600000 336.350000 ;
      RECT 0.000000 335.550000 697.600000 336.050000 ;
      RECT 0.720000 335.250000 697.600000 335.550000 ;
      RECT 0.000000 334.750000 697.600000 335.250000 ;
      RECT 0.720000 334.450000 697.600000 334.750000 ;
      RECT 0.000000 333.950000 697.600000 334.450000 ;
      RECT 0.720000 333.650000 697.600000 333.950000 ;
      RECT 0.000000 333.150000 697.600000 333.650000 ;
      RECT 0.720000 332.850000 697.600000 333.150000 ;
      RECT 0.000000 332.350000 697.600000 332.850000 ;
      RECT 0.720000 332.050000 697.600000 332.350000 ;
      RECT 0.000000 331.550000 697.600000 332.050000 ;
      RECT 0.720000 331.250000 697.600000 331.550000 ;
      RECT 0.000000 330.750000 697.600000 331.250000 ;
      RECT 0.720000 330.450000 697.600000 330.750000 ;
      RECT 0.000000 329.950000 697.600000 330.450000 ;
      RECT 0.720000 329.650000 697.600000 329.950000 ;
      RECT 0.000000 329.150000 697.600000 329.650000 ;
      RECT 0.720000 328.850000 697.600000 329.150000 ;
      RECT 0.000000 328.350000 697.600000 328.850000 ;
      RECT 0.720000 328.050000 697.600000 328.350000 ;
      RECT 0.000000 327.550000 697.600000 328.050000 ;
      RECT 0.720000 327.250000 697.600000 327.550000 ;
      RECT 0.000000 326.750000 697.600000 327.250000 ;
      RECT 0.720000 326.450000 697.600000 326.750000 ;
      RECT 0.000000 325.950000 697.600000 326.450000 ;
      RECT 0.720000 325.650000 697.600000 325.950000 ;
      RECT 0.000000 325.150000 697.600000 325.650000 ;
      RECT 0.720000 324.850000 697.600000 325.150000 ;
      RECT 0.000000 324.350000 697.600000 324.850000 ;
      RECT 0.720000 324.050000 697.600000 324.350000 ;
      RECT 0.000000 323.550000 697.600000 324.050000 ;
      RECT 0.720000 323.250000 697.600000 323.550000 ;
      RECT 0.000000 322.750000 697.600000 323.250000 ;
      RECT 0.720000 322.450000 697.600000 322.750000 ;
      RECT 0.000000 321.950000 697.600000 322.450000 ;
      RECT 0.720000 321.650000 697.600000 321.950000 ;
      RECT 0.000000 321.150000 697.600000 321.650000 ;
      RECT 0.720000 320.850000 697.600000 321.150000 ;
      RECT 0.000000 320.350000 697.600000 320.850000 ;
      RECT 0.720000 320.050000 697.600000 320.350000 ;
      RECT 0.000000 319.550000 697.600000 320.050000 ;
      RECT 0.720000 319.250000 697.600000 319.550000 ;
      RECT 0.000000 318.750000 697.600000 319.250000 ;
      RECT 0.720000 318.450000 697.600000 318.750000 ;
      RECT 0.000000 317.950000 697.600000 318.450000 ;
      RECT 0.720000 317.650000 697.600000 317.950000 ;
      RECT 0.000000 317.150000 697.600000 317.650000 ;
      RECT 0.720000 316.850000 697.600000 317.150000 ;
      RECT 0.000000 316.350000 697.600000 316.850000 ;
      RECT 0.720000 316.050000 697.600000 316.350000 ;
      RECT 0.000000 315.550000 697.600000 316.050000 ;
      RECT 0.720000 315.250000 697.600000 315.550000 ;
      RECT 0.000000 314.750000 697.600000 315.250000 ;
      RECT 0.720000 314.450000 697.600000 314.750000 ;
      RECT 0.000000 313.950000 697.600000 314.450000 ;
      RECT 0.720000 313.650000 697.600000 313.950000 ;
      RECT 0.000000 313.150000 697.600000 313.650000 ;
      RECT 0.720000 312.850000 697.600000 313.150000 ;
      RECT 0.000000 312.350000 697.600000 312.850000 ;
      RECT 0.720000 312.050000 697.600000 312.350000 ;
      RECT 0.000000 311.550000 697.600000 312.050000 ;
      RECT 0.720000 311.250000 697.600000 311.550000 ;
      RECT 0.000000 310.750000 697.600000 311.250000 ;
      RECT 0.720000 310.450000 697.600000 310.750000 ;
      RECT 0.000000 309.950000 697.600000 310.450000 ;
      RECT 0.720000 309.650000 697.600000 309.950000 ;
      RECT 0.000000 309.150000 697.600000 309.650000 ;
      RECT 0.720000 308.850000 697.600000 309.150000 ;
      RECT 0.000000 308.350000 697.600000 308.850000 ;
      RECT 0.720000 308.050000 697.600000 308.350000 ;
      RECT 0.000000 307.550000 697.600000 308.050000 ;
      RECT 0.720000 307.250000 697.600000 307.550000 ;
      RECT 0.000000 306.750000 697.600000 307.250000 ;
      RECT 0.720000 306.450000 697.600000 306.750000 ;
      RECT 0.000000 305.950000 697.600000 306.450000 ;
      RECT 0.720000 305.650000 697.600000 305.950000 ;
      RECT 0.000000 305.150000 697.600000 305.650000 ;
      RECT 0.720000 304.850000 697.600000 305.150000 ;
      RECT 0.000000 304.350000 697.600000 304.850000 ;
      RECT 0.720000 304.050000 697.600000 304.350000 ;
      RECT 0.000000 303.550000 697.600000 304.050000 ;
      RECT 0.720000 303.250000 697.600000 303.550000 ;
      RECT 0.000000 302.750000 697.600000 303.250000 ;
      RECT 0.720000 302.450000 697.600000 302.750000 ;
      RECT 0.000000 301.950000 697.600000 302.450000 ;
      RECT 0.720000 301.650000 697.600000 301.950000 ;
      RECT 0.000000 301.150000 697.600000 301.650000 ;
      RECT 0.720000 300.850000 697.600000 301.150000 ;
      RECT 0.000000 300.350000 697.600000 300.850000 ;
      RECT 0.720000 300.050000 697.600000 300.350000 ;
      RECT 0.000000 299.550000 697.600000 300.050000 ;
      RECT 0.720000 299.250000 697.600000 299.550000 ;
      RECT 0.000000 298.750000 697.600000 299.250000 ;
      RECT 0.720000 298.450000 697.600000 298.750000 ;
      RECT 0.000000 297.950000 697.600000 298.450000 ;
      RECT 0.720000 297.650000 697.600000 297.950000 ;
      RECT 0.000000 297.150000 697.600000 297.650000 ;
      RECT 0.720000 296.850000 697.600000 297.150000 ;
      RECT 0.000000 296.350000 697.600000 296.850000 ;
      RECT 0.720000 296.050000 697.600000 296.350000 ;
      RECT 0.000000 295.550000 697.600000 296.050000 ;
      RECT 0.720000 295.250000 697.600000 295.550000 ;
      RECT 0.000000 294.750000 697.600000 295.250000 ;
      RECT 0.720000 294.450000 697.600000 294.750000 ;
      RECT 0.000000 293.950000 697.600000 294.450000 ;
      RECT 0.720000 293.650000 697.600000 293.950000 ;
      RECT 0.000000 293.150000 697.600000 293.650000 ;
      RECT 0.720000 292.850000 697.600000 293.150000 ;
      RECT 0.000000 292.350000 697.600000 292.850000 ;
      RECT 0.720000 292.050000 697.600000 292.350000 ;
      RECT 0.000000 291.550000 697.600000 292.050000 ;
      RECT 0.720000 291.250000 697.600000 291.550000 ;
      RECT 0.000000 290.750000 697.600000 291.250000 ;
      RECT 0.720000 290.450000 697.600000 290.750000 ;
      RECT 0.000000 289.950000 697.600000 290.450000 ;
      RECT 0.720000 289.650000 697.600000 289.950000 ;
      RECT 0.000000 289.150000 697.600000 289.650000 ;
      RECT 0.720000 288.850000 697.600000 289.150000 ;
      RECT 0.000000 0.760000 697.600000 288.850000 ;
      RECT 422.310000 0.000000 697.600000 0.760000 ;
      RECT 421.510000 0.000000 421.890000 0.760000 ;
      RECT 420.710000 0.000000 421.090000 0.760000 ;
      RECT 419.910000 0.000000 420.290000 0.760000 ;
      RECT 419.110000 0.000000 419.490000 0.760000 ;
      RECT 418.310000 0.000000 418.690000 0.760000 ;
      RECT 417.510000 0.000000 417.890000 0.760000 ;
      RECT 416.710000 0.000000 417.090000 0.760000 ;
      RECT 415.910000 0.000000 416.290000 0.760000 ;
      RECT 415.110000 0.000000 415.490000 0.760000 ;
      RECT 414.310000 0.000000 414.690000 0.760000 ;
      RECT 413.510000 0.000000 413.890000 0.760000 ;
      RECT 412.710000 0.000000 413.090000 0.760000 ;
      RECT 411.910000 0.000000 412.290000 0.760000 ;
      RECT 411.110000 0.000000 411.490000 0.760000 ;
      RECT 410.310000 0.000000 410.690000 0.760000 ;
      RECT 409.510000 0.000000 409.890000 0.760000 ;
      RECT 408.710000 0.000000 409.090000 0.760000 ;
      RECT 407.910000 0.000000 408.290000 0.760000 ;
      RECT 407.110000 0.000000 407.490000 0.760000 ;
      RECT 406.310000 0.000000 406.690000 0.760000 ;
      RECT 405.510000 0.000000 405.890000 0.760000 ;
      RECT 404.710000 0.000000 405.090000 0.760000 ;
      RECT 403.910000 0.000000 404.290000 0.760000 ;
      RECT 403.110000 0.000000 403.490000 0.760000 ;
      RECT 402.310000 0.000000 402.690000 0.760000 ;
      RECT 401.510000 0.000000 401.890000 0.760000 ;
      RECT 400.710000 0.000000 401.090000 0.760000 ;
      RECT 399.910000 0.000000 400.290000 0.760000 ;
      RECT 399.110000 0.000000 399.490000 0.760000 ;
      RECT 398.310000 0.000000 398.690000 0.760000 ;
      RECT 397.510000 0.000000 397.890000 0.760000 ;
      RECT 396.710000 0.000000 397.090000 0.760000 ;
      RECT 395.910000 0.000000 396.290000 0.760000 ;
      RECT 395.110000 0.000000 395.490000 0.760000 ;
      RECT 394.310000 0.000000 394.690000 0.760000 ;
      RECT 393.510000 0.000000 393.890000 0.760000 ;
      RECT 392.710000 0.000000 393.090000 0.760000 ;
      RECT 391.910000 0.000000 392.290000 0.760000 ;
      RECT 391.110000 0.000000 391.490000 0.760000 ;
      RECT 390.310000 0.000000 390.690000 0.760000 ;
      RECT 389.510000 0.000000 389.890000 0.760000 ;
      RECT 388.710000 0.000000 389.090000 0.760000 ;
      RECT 387.910000 0.000000 388.290000 0.760000 ;
      RECT 387.110000 0.000000 387.490000 0.760000 ;
      RECT 386.310000 0.000000 386.690000 0.760000 ;
      RECT 385.510000 0.000000 385.890000 0.760000 ;
      RECT 384.710000 0.000000 385.090000 0.760000 ;
      RECT 383.910000 0.000000 384.290000 0.760000 ;
      RECT 383.110000 0.000000 383.490000 0.760000 ;
      RECT 382.310000 0.000000 382.690000 0.760000 ;
      RECT 381.510000 0.000000 381.890000 0.760000 ;
      RECT 380.710000 0.000000 381.090000 0.760000 ;
      RECT 379.910000 0.000000 380.290000 0.760000 ;
      RECT 379.110000 0.000000 379.490000 0.760000 ;
      RECT 378.310000 0.000000 378.690000 0.760000 ;
      RECT 377.510000 0.000000 377.890000 0.760000 ;
      RECT 376.710000 0.000000 377.090000 0.760000 ;
      RECT 375.910000 0.000000 376.290000 0.760000 ;
      RECT 375.110000 0.000000 375.490000 0.760000 ;
      RECT 374.310000 0.000000 374.690000 0.760000 ;
      RECT 373.510000 0.000000 373.890000 0.760000 ;
      RECT 372.710000 0.000000 373.090000 0.760000 ;
      RECT 371.910000 0.000000 372.290000 0.760000 ;
      RECT 371.110000 0.000000 371.490000 0.760000 ;
      RECT 370.310000 0.000000 370.690000 0.760000 ;
      RECT 369.510000 0.000000 369.890000 0.760000 ;
      RECT 368.710000 0.000000 369.090000 0.760000 ;
      RECT 367.910000 0.000000 368.290000 0.760000 ;
      RECT 367.110000 0.000000 367.490000 0.760000 ;
      RECT 366.310000 0.000000 366.690000 0.760000 ;
      RECT 365.510000 0.000000 365.890000 0.760000 ;
      RECT 364.710000 0.000000 365.090000 0.760000 ;
      RECT 363.910000 0.000000 364.290000 0.760000 ;
      RECT 363.110000 0.000000 363.490000 0.760000 ;
      RECT 362.310000 0.000000 362.690000 0.760000 ;
      RECT 361.510000 0.000000 361.890000 0.760000 ;
      RECT 360.710000 0.000000 361.090000 0.760000 ;
      RECT 359.910000 0.000000 360.290000 0.760000 ;
      RECT 359.110000 0.000000 359.490000 0.760000 ;
      RECT 358.310000 0.000000 358.690000 0.760000 ;
      RECT 357.510000 0.000000 357.890000 0.760000 ;
      RECT 356.710000 0.000000 357.090000 0.760000 ;
      RECT 355.910000 0.000000 356.290000 0.760000 ;
      RECT 355.110000 0.000000 355.490000 0.760000 ;
      RECT 354.310000 0.000000 354.690000 0.760000 ;
      RECT 353.510000 0.000000 353.890000 0.760000 ;
      RECT 352.710000 0.000000 353.090000 0.760000 ;
      RECT 351.910000 0.000000 352.290000 0.760000 ;
      RECT 351.110000 0.000000 351.490000 0.760000 ;
      RECT 350.310000 0.000000 350.690000 0.760000 ;
      RECT 349.510000 0.000000 349.890000 0.760000 ;
      RECT 348.710000 0.000000 349.090000 0.760000 ;
      RECT 347.910000 0.000000 348.290000 0.760000 ;
      RECT 347.110000 0.000000 347.490000 0.760000 ;
      RECT 346.310000 0.000000 346.690000 0.760000 ;
      RECT 345.510000 0.000000 345.890000 0.760000 ;
      RECT 344.710000 0.000000 345.090000 0.760000 ;
      RECT 343.910000 0.000000 344.290000 0.760000 ;
      RECT 343.110000 0.000000 343.490000 0.760000 ;
      RECT 342.310000 0.000000 342.690000 0.760000 ;
      RECT 341.510000 0.000000 341.890000 0.760000 ;
      RECT 340.710000 0.000000 341.090000 0.760000 ;
      RECT 339.910000 0.000000 340.290000 0.760000 ;
      RECT 339.110000 0.000000 339.490000 0.760000 ;
      RECT 338.310000 0.000000 338.690000 0.760000 ;
      RECT 337.510000 0.000000 337.890000 0.760000 ;
      RECT 336.710000 0.000000 337.090000 0.760000 ;
      RECT 335.910000 0.000000 336.290000 0.760000 ;
      RECT 335.110000 0.000000 335.490000 0.760000 ;
      RECT 334.310000 0.000000 334.690000 0.760000 ;
      RECT 333.510000 0.000000 333.890000 0.760000 ;
      RECT 332.710000 0.000000 333.090000 0.760000 ;
      RECT 331.910000 0.000000 332.290000 0.760000 ;
      RECT 331.110000 0.000000 331.490000 0.760000 ;
      RECT 330.310000 0.000000 330.690000 0.760000 ;
      RECT 329.510000 0.000000 329.890000 0.760000 ;
      RECT 328.710000 0.000000 329.090000 0.760000 ;
      RECT 327.910000 0.000000 328.290000 0.760000 ;
      RECT 327.110000 0.000000 327.490000 0.760000 ;
      RECT 326.310000 0.000000 326.690000 0.760000 ;
      RECT 325.510000 0.000000 325.890000 0.760000 ;
      RECT 324.710000 0.000000 325.090000 0.760000 ;
      RECT 323.910000 0.000000 324.290000 0.760000 ;
      RECT 323.110000 0.000000 323.490000 0.760000 ;
      RECT 322.310000 0.000000 322.690000 0.760000 ;
      RECT 321.510000 0.000000 321.890000 0.760000 ;
      RECT 320.710000 0.000000 321.090000 0.760000 ;
      RECT 319.910000 0.000000 320.290000 0.760000 ;
      RECT 319.110000 0.000000 319.490000 0.760000 ;
      RECT 318.310000 0.000000 318.690000 0.760000 ;
      RECT 317.510000 0.000000 317.890000 0.760000 ;
      RECT 316.710000 0.000000 317.090000 0.760000 ;
      RECT 315.910000 0.000000 316.290000 0.760000 ;
      RECT 315.110000 0.000000 315.490000 0.760000 ;
      RECT 314.310000 0.000000 314.690000 0.760000 ;
      RECT 313.510000 0.000000 313.890000 0.760000 ;
      RECT 312.710000 0.000000 313.090000 0.760000 ;
      RECT 311.910000 0.000000 312.290000 0.760000 ;
      RECT 311.110000 0.000000 311.490000 0.760000 ;
      RECT 310.310000 0.000000 310.690000 0.760000 ;
      RECT 309.510000 0.000000 309.890000 0.760000 ;
      RECT 308.710000 0.000000 309.090000 0.760000 ;
      RECT 307.910000 0.000000 308.290000 0.760000 ;
      RECT 307.110000 0.000000 307.490000 0.760000 ;
      RECT 306.310000 0.000000 306.690000 0.760000 ;
      RECT 305.510000 0.000000 305.890000 0.760000 ;
      RECT 304.710000 0.000000 305.090000 0.760000 ;
      RECT 303.910000 0.000000 304.290000 0.760000 ;
      RECT 303.110000 0.000000 303.490000 0.760000 ;
      RECT 302.310000 0.000000 302.690000 0.760000 ;
      RECT 301.510000 0.000000 301.890000 0.760000 ;
      RECT 300.710000 0.000000 301.090000 0.760000 ;
      RECT 299.910000 0.000000 300.290000 0.760000 ;
      RECT 299.110000 0.000000 299.490000 0.760000 ;
      RECT 298.310000 0.000000 298.690000 0.760000 ;
      RECT 297.510000 0.000000 297.890000 0.760000 ;
      RECT 296.710000 0.000000 297.090000 0.760000 ;
      RECT 295.910000 0.000000 296.290000 0.760000 ;
      RECT 295.110000 0.000000 295.490000 0.760000 ;
      RECT 294.310000 0.000000 294.690000 0.760000 ;
      RECT 293.510000 0.000000 293.890000 0.760000 ;
      RECT 292.710000 0.000000 293.090000 0.760000 ;
      RECT 291.910000 0.000000 292.290000 0.760000 ;
      RECT 291.110000 0.000000 291.490000 0.760000 ;
      RECT 290.310000 0.000000 290.690000 0.760000 ;
      RECT 289.510000 0.000000 289.890000 0.760000 ;
      RECT 288.710000 0.000000 289.090000 0.760000 ;
      RECT 287.910000 0.000000 288.290000 0.760000 ;
      RECT 287.110000 0.000000 287.490000 0.760000 ;
      RECT 286.310000 0.000000 286.690000 0.760000 ;
      RECT 285.510000 0.000000 285.890000 0.760000 ;
      RECT 284.710000 0.000000 285.090000 0.760000 ;
      RECT 283.910000 0.000000 284.290000 0.760000 ;
      RECT 283.110000 0.000000 283.490000 0.760000 ;
      RECT 282.310000 0.000000 282.690000 0.760000 ;
      RECT 281.510000 0.000000 281.890000 0.760000 ;
      RECT 280.710000 0.000000 281.090000 0.760000 ;
      RECT 279.910000 0.000000 280.290000 0.760000 ;
      RECT 279.110000 0.000000 279.490000 0.760000 ;
      RECT 278.310000 0.000000 278.690000 0.760000 ;
      RECT 277.510000 0.000000 277.890000 0.760000 ;
      RECT 276.710000 0.000000 277.090000 0.760000 ;
      RECT 275.910000 0.000000 276.290000 0.760000 ;
      RECT 0.000000 0.000000 275.490000 0.760000 ;
    LAYER M4 ;
      RECT 0.000000 0.000000 697.600000 695.000000 ;
    LAYER M5 ;
      RECT 0.000000 0.000000 697.600000 695.000000 ;
    LAYER M6 ;
      RECT 0.000000 0.000000 697.600000 695.000000 ;
    LAYER M7 ;
      RECT 0.000000 0.000000 697.600000 695.000000 ;
    LAYER M8 ;
      RECT 0.000000 0.000000 697.600000 695.000000 ;
  END
END fullchip

END LIBRARY
