##
## LEF for PtnCells ;
## created by Innovus v19.17-s077_1 on Sat Mar 18 23:18:39 2023
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO fullchip
  CLASS BLOCK ;
  SIZE 394.600000 BY 394.400000 ;
  FOREIGN fullchip 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 150.950000 0.600000 151.050000 ;
    END
  END clk
  PIN mem_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 241.950000 0.600000 242.050000 ;
    END
  END mem_in[63]
  PIN mem_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 240.950000 0.600000 241.050000 ;
    END
  END mem_in[62]
  PIN mem_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 239.950000 0.600000 240.050000 ;
    END
  END mem_in[61]
  PIN mem_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 238.950000 0.600000 239.050000 ;
    END
  END mem_in[60]
  PIN mem_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 237.950000 0.600000 238.050000 ;
    END
  END mem_in[59]
  PIN mem_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 236.950000 0.600000 237.050000 ;
    END
  END mem_in[58]
  PIN mem_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 235.950000 0.600000 236.050000 ;
    END
  END mem_in[57]
  PIN mem_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 234.950000 0.600000 235.050000 ;
    END
  END mem_in[56]
  PIN mem_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 233.950000 0.600000 234.050000 ;
    END
  END mem_in[55]
  PIN mem_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 232.950000 0.600000 233.050000 ;
    END
  END mem_in[54]
  PIN mem_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 231.950000 0.600000 232.050000 ;
    END
  END mem_in[53]
  PIN mem_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 230.950000 0.600000 231.050000 ;
    END
  END mem_in[52]
  PIN mem_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 229.950000 0.600000 230.050000 ;
    END
  END mem_in[51]
  PIN mem_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 228.950000 0.600000 229.050000 ;
    END
  END mem_in[50]
  PIN mem_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 227.950000 0.600000 228.050000 ;
    END
  END mem_in[49]
  PIN mem_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 226.950000 0.600000 227.050000 ;
    END
  END mem_in[48]
  PIN mem_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 225.950000 0.600000 226.050000 ;
    END
  END mem_in[47]
  PIN mem_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 224.950000 0.600000 225.050000 ;
    END
  END mem_in[46]
  PIN mem_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 223.950000 0.600000 224.050000 ;
    END
  END mem_in[45]
  PIN mem_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 222.950000 0.600000 223.050000 ;
    END
  END mem_in[44]
  PIN mem_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 221.950000 0.600000 222.050000 ;
    END
  END mem_in[43]
  PIN mem_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 220.950000 0.600000 221.050000 ;
    END
  END mem_in[42]
  PIN mem_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 219.950000 0.600000 220.050000 ;
    END
  END mem_in[41]
  PIN mem_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 218.950000 0.600000 219.050000 ;
    END
  END mem_in[40]
  PIN mem_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 217.950000 0.600000 218.050000 ;
    END
  END mem_in[39]
  PIN mem_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 216.950000 0.600000 217.050000 ;
    END
  END mem_in[38]
  PIN mem_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 215.950000 0.600000 216.050000 ;
    END
  END mem_in[37]
  PIN mem_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 214.950000 0.600000 215.050000 ;
    END
  END mem_in[36]
  PIN mem_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 213.950000 0.600000 214.050000 ;
    END
  END mem_in[35]
  PIN mem_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 212.950000 0.600000 213.050000 ;
    END
  END mem_in[34]
  PIN mem_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 211.950000 0.600000 212.050000 ;
    END
  END mem_in[33]
  PIN mem_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 210.950000 0.600000 211.050000 ;
    END
  END mem_in[32]
  PIN mem_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 209.950000 0.600000 210.050000 ;
    END
  END mem_in[31]
  PIN mem_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 208.950000 0.600000 209.050000 ;
    END
  END mem_in[30]
  PIN mem_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 207.950000 0.600000 208.050000 ;
    END
  END mem_in[29]
  PIN mem_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 206.950000 0.600000 207.050000 ;
    END
  END mem_in[28]
  PIN mem_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 205.950000 0.600000 206.050000 ;
    END
  END mem_in[27]
  PIN mem_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 204.950000 0.600000 205.050000 ;
    END
  END mem_in[26]
  PIN mem_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 203.950000 0.600000 204.050000 ;
    END
  END mem_in[25]
  PIN mem_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 202.950000 0.600000 203.050000 ;
    END
  END mem_in[24]
  PIN mem_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 201.950000 0.600000 202.050000 ;
    END
  END mem_in[23]
  PIN mem_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 200.950000 0.600000 201.050000 ;
    END
  END mem_in[22]
  PIN mem_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 199.950000 0.600000 200.050000 ;
    END
  END mem_in[21]
  PIN mem_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 198.950000 0.600000 199.050000 ;
    END
  END mem_in[20]
  PIN mem_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 197.950000 0.600000 198.050000 ;
    END
  END mem_in[19]
  PIN mem_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 196.950000 0.600000 197.050000 ;
    END
  END mem_in[18]
  PIN mem_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 195.950000 0.600000 196.050000 ;
    END
  END mem_in[17]
  PIN mem_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 194.950000 0.600000 195.050000 ;
    END
  END mem_in[16]
  PIN mem_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 193.950000 0.600000 194.050000 ;
    END
  END mem_in[15]
  PIN mem_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 192.950000 0.600000 193.050000 ;
    END
  END mem_in[14]
  PIN mem_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 191.950000 0.600000 192.050000 ;
    END
  END mem_in[13]
  PIN mem_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 190.950000 0.600000 191.050000 ;
    END
  END mem_in[12]
  PIN mem_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 189.950000 0.600000 190.050000 ;
    END
  END mem_in[11]
  PIN mem_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 188.950000 0.600000 189.050000 ;
    END
  END mem_in[10]
  PIN mem_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 187.950000 0.600000 188.050000 ;
    END
  END mem_in[9]
  PIN mem_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 186.950000 0.600000 187.050000 ;
    END
  END mem_in[8]
  PIN mem_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 185.950000 0.600000 186.050000 ;
    END
  END mem_in[7]
  PIN mem_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 184.950000 0.600000 185.050000 ;
    END
  END mem_in[6]
  PIN mem_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 183.950000 0.600000 184.050000 ;
    END
  END mem_in[5]
  PIN mem_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 182.950000 0.600000 183.050000 ;
    END
  END mem_in[4]
  PIN mem_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 181.950000 0.600000 182.050000 ;
    END
  END mem_in[3]
  PIN mem_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 180.950000 0.600000 181.050000 ;
    END
  END mem_in[2]
  PIN mem_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 179.950000 0.600000 180.050000 ;
    END
  END mem_in[1]
  PIN mem_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 178.950000 0.600000 179.050000 ;
    END
  END mem_in[0]
  PIN inst[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 177.950000 0.600000 178.050000 ;
    END
  END inst[26]
  PIN inst[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 176.950000 0.600000 177.050000 ;
    END
  END inst[25]
  PIN inst[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 175.950000 0.600000 176.050000 ;
    END
  END inst[24]
  PIN inst[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 174.950000 0.600000 175.050000 ;
    END
  END inst[23]
  PIN inst[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 173.950000 0.600000 174.050000 ;
    END
  END inst[22]
  PIN inst[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 172.950000 0.600000 173.050000 ;
    END
  END inst[21]
  PIN inst[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 171.950000 0.600000 172.050000 ;
    END
  END inst[20]
  PIN inst[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 170.950000 0.600000 171.050000 ;
    END
  END inst[19]
  PIN inst[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 169.950000 0.600000 170.050000 ;
    END
  END inst[18]
  PIN inst[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 168.950000 0.600000 169.050000 ;
    END
  END inst[17]
  PIN inst[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 167.950000 0.600000 168.050000 ;
    END
  END inst[16]
  PIN inst[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 166.950000 0.600000 167.050000 ;
    END
  END inst[15]
  PIN inst[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 165.950000 0.600000 166.050000 ;
    END
  END inst[14]
  PIN inst[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 164.950000 0.600000 165.050000 ;
    END
  END inst[13]
  PIN inst[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 163.950000 0.600000 164.050000 ;
    END
  END inst[12]
  PIN inst[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 162.950000 0.600000 163.050000 ;
    END
  END inst[11]
  PIN inst[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 161.950000 0.600000 162.050000 ;
    END
  END inst[10]
  PIN inst[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 160.950000 0.600000 161.050000 ;
    END
  END inst[9]
  PIN inst[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 159.950000 0.600000 160.050000 ;
    END
  END inst[8]
  PIN inst[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 158.950000 0.600000 159.050000 ;
    END
  END inst[7]
  PIN inst[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 157.950000 0.600000 158.050000 ;
    END
  END inst[6]
  PIN inst[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 156.950000 0.600000 157.050000 ;
    END
  END inst[5]
  PIN inst[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 155.950000 0.600000 156.050000 ;
    END
  END inst[4]
  PIN inst[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 154.950000 0.600000 155.050000 ;
    END
  END inst[3]
  PIN inst[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 153.950000 0.600000 154.050000 ;
    END
  END inst[2]
  PIN inst[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 152.950000 0.600000 153.050000 ;
    END
  END inst[1]
  PIN inst[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 151.950000 0.600000 152.050000 ;
    END
  END inst[0]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.000000 242.950000 0.600000 243.050000 ;
    END
  END reset
  PIN out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 236.450000 0.000000 236.550000 0.600000 ;
    END
  END out[95]
  PIN out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 235.450000 0.000000 235.550000 0.600000 ;
    END
  END out[94]
  PIN out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 234.450000 0.000000 234.550000 0.600000 ;
    END
  END out[93]
  PIN out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 233.450000 0.000000 233.550000 0.600000 ;
    END
  END out[92]
  PIN out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 232.450000 0.000000 232.550000 0.600000 ;
    END
  END out[91]
  PIN out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 231.450000 0.000000 231.550000 0.600000 ;
    END
  END out[90]
  PIN out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 230.450000 0.000000 230.550000 0.600000 ;
    END
  END out[89]
  PIN out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 229.450000 0.000000 229.550000 0.600000 ;
    END
  END out[88]
  PIN out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 228.450000 0.000000 228.550000 0.600000 ;
    END
  END out[87]
  PIN out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 227.450000 0.000000 227.550000 0.600000 ;
    END
  END out[86]
  PIN out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 226.450000 0.000000 226.550000 0.600000 ;
    END
  END out[85]
  PIN out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 225.450000 0.000000 225.550000 0.600000 ;
    END
  END out[84]
  PIN out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 224.450000 0.000000 224.550000 0.600000 ;
    END
  END out[83]
  PIN out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 223.450000 0.000000 223.550000 0.600000 ;
    END
  END out[82]
  PIN out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 222.450000 0.000000 222.550000 0.600000 ;
    END
  END out[81]
  PIN out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 221.450000 0.000000 221.550000 0.600000 ;
    END
  END out[80]
  PIN out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 220.450000 0.000000 220.550000 0.600000 ;
    END
  END out[79]
  PIN out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 219.450000 0.000000 219.550000 0.600000 ;
    END
  END out[78]
  PIN out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 218.450000 0.000000 218.550000 0.600000 ;
    END
  END out[77]
  PIN out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 217.450000 0.000000 217.550000 0.600000 ;
    END
  END out[76]
  PIN out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 216.450000 0.000000 216.550000 0.600000 ;
    END
  END out[75]
  PIN out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 215.450000 0.000000 215.550000 0.600000 ;
    END
  END out[74]
  PIN out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 214.450000 0.000000 214.550000 0.600000 ;
    END
  END out[73]
  PIN out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 213.450000 0.000000 213.550000 0.600000 ;
    END
  END out[72]
  PIN out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 212.450000 0.000000 212.550000 0.600000 ;
    END
  END out[71]
  PIN out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 211.450000 0.000000 211.550000 0.600000 ;
    END
  END out[70]
  PIN out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 210.450000 0.000000 210.550000 0.600000 ;
    END
  END out[69]
  PIN out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 209.450000 0.000000 209.550000 0.600000 ;
    END
  END out[68]
  PIN out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 208.450000 0.000000 208.550000 0.600000 ;
    END
  END out[67]
  PIN out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 207.450000 0.000000 207.550000 0.600000 ;
    END
  END out[66]
  PIN out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 206.450000 0.000000 206.550000 0.600000 ;
    END
  END out[65]
  PIN out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 205.450000 0.000000 205.550000 0.600000 ;
    END
  END out[64]
  PIN out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 204.450000 0.000000 204.550000 0.600000 ;
    END
  END out[63]
  PIN out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 203.450000 0.000000 203.550000 0.600000 ;
    END
  END out[62]
  PIN out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 202.450000 0.000000 202.550000 0.600000 ;
    END
  END out[61]
  PIN out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 201.450000 0.000000 201.550000 0.600000 ;
    END
  END out[60]
  PIN out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 200.450000 0.000000 200.550000 0.600000 ;
    END
  END out[59]
  PIN out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 199.450000 0.000000 199.550000 0.600000 ;
    END
  END out[58]
  PIN out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 198.450000 0.000000 198.550000 0.600000 ;
    END
  END out[57]
  PIN out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 197.450000 0.000000 197.550000 0.600000 ;
    END
  END out[56]
  PIN out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 196.450000 0.000000 196.550000 0.600000 ;
    END
  END out[55]
  PIN out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 195.450000 0.000000 195.550000 0.600000 ;
    END
  END out[54]
  PIN out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 194.450000 0.000000 194.550000 0.600000 ;
    END
  END out[53]
  PIN out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 193.450000 0.000000 193.550000 0.600000 ;
    END
  END out[52]
  PIN out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 192.450000 0.000000 192.550000 0.600000 ;
    END
  END out[51]
  PIN out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 191.450000 0.000000 191.550000 0.600000 ;
    END
  END out[50]
  PIN out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 190.450000 0.000000 190.550000 0.600000 ;
    END
  END out[49]
  PIN out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 189.450000 0.000000 189.550000 0.600000 ;
    END
  END out[48]
  PIN out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 188.450000 0.000000 188.550000 0.600000 ;
    END
  END out[47]
  PIN out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 187.450000 0.000000 187.550000 0.600000 ;
    END
  END out[46]
  PIN out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 186.450000 0.000000 186.550000 0.600000 ;
    END
  END out[45]
  PIN out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 185.450000 0.000000 185.550000 0.600000 ;
    END
  END out[44]
  PIN out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 184.450000 0.000000 184.550000 0.600000 ;
    END
  END out[43]
  PIN out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 183.450000 0.000000 183.550000 0.600000 ;
    END
  END out[42]
  PIN out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 182.450000 0.000000 182.550000 0.600000 ;
    END
  END out[41]
  PIN out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 181.450000 0.000000 181.550000 0.600000 ;
    END
  END out[40]
  PIN out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 180.450000 0.000000 180.550000 0.600000 ;
    END
  END out[39]
  PIN out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 179.450000 0.000000 179.550000 0.600000 ;
    END
  END out[38]
  PIN out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 178.450000 0.000000 178.550000 0.600000 ;
    END
  END out[37]
  PIN out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 177.450000 0.000000 177.550000 0.600000 ;
    END
  END out[36]
  PIN out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 176.450000 0.000000 176.550000 0.600000 ;
    END
  END out[35]
  PIN out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 175.450000 0.000000 175.550000 0.600000 ;
    END
  END out[34]
  PIN out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 174.450000 0.000000 174.550000 0.600000 ;
    END
  END out[33]
  PIN out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 173.450000 0.000000 173.550000 0.600000 ;
    END
  END out[32]
  PIN out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 172.450000 0.000000 172.550000 0.600000 ;
    END
  END out[31]
  PIN out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 171.450000 0.000000 171.550000 0.600000 ;
    END
  END out[30]
  PIN out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 170.450000 0.000000 170.550000 0.600000 ;
    END
  END out[29]
  PIN out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 169.450000 0.000000 169.550000 0.600000 ;
    END
  END out[28]
  PIN out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 168.450000 0.000000 168.550000 0.600000 ;
    END
  END out[27]
  PIN out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 167.450000 0.000000 167.550000 0.600000 ;
    END
  END out[26]
  PIN out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 166.450000 0.000000 166.550000 0.600000 ;
    END
  END out[25]
  PIN out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 165.450000 0.000000 165.550000 0.600000 ;
    END
  END out[24]
  PIN out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 164.450000 0.000000 164.550000 0.600000 ;
    END
  END out[23]
  PIN out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 163.450000 0.000000 163.550000 0.600000 ;
    END
  END out[22]
  PIN out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 162.450000 0.000000 162.550000 0.600000 ;
    END
  END out[21]
  PIN out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 161.450000 0.000000 161.550000 0.600000 ;
    END
  END out[20]
  PIN out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 160.450000 0.000000 160.550000 0.600000 ;
    END
  END out[19]
  PIN out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 159.450000 0.000000 159.550000 0.600000 ;
    END
  END out[18]
  PIN out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 158.450000 0.000000 158.550000 0.600000 ;
    END
  END out[17]
  PIN out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 157.450000 0.000000 157.550000 0.600000 ;
    END
  END out[16]
  PIN out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 156.450000 0.000000 156.550000 0.600000 ;
    END
  END out[15]
  PIN out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 155.450000 0.000000 155.550000 0.600000 ;
    END
  END out[14]
  PIN out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 154.450000 0.000000 154.550000 0.600000 ;
    END
  END out[13]
  PIN out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 153.450000 0.000000 153.550000 0.600000 ;
    END
  END out[12]
  PIN out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 152.450000 0.000000 152.550000 0.600000 ;
    END
  END out[11]
  PIN out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 151.450000 0.000000 151.550000 0.600000 ;
    END
  END out[10]
  PIN out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 150.450000 0.000000 150.550000 0.600000 ;
    END
  END out[9]
  PIN out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 149.450000 0.000000 149.550000 0.600000 ;
    END
  END out[8]
  PIN out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 148.450000 0.000000 148.550000 0.600000 ;
    END
  END out[7]
  PIN out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 147.450000 0.000000 147.550000 0.600000 ;
    END
  END out[6]
  PIN out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 146.450000 0.000000 146.550000 0.600000 ;
    END
  END out[5]
  PIN out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 145.450000 0.000000 145.550000 0.600000 ;
    END
  END out[4]
  PIN out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 144.450000 0.000000 144.550000 0.600000 ;
    END
  END out[3]
  PIN out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 143.450000 0.000000 143.550000 0.600000 ;
    END
  END out[2]
  PIN out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 142.450000 0.000000 142.550000 0.600000 ;
    END
  END out[1]
  PIN out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 141.450000 0.000000 141.550000 0.600000 ;
    END
  END out[0]
  PIN sum_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 252.450000 0.000000 252.550000 0.600000 ;
    END
  END sum_out[15]
  PIN sum_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 251.450000 0.000000 251.550000 0.600000 ;
    END
  END sum_out[14]
  PIN sum_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 250.450000 0.000000 250.550000 0.600000 ;
    END
  END sum_out[13]
  PIN sum_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 249.450000 0.000000 249.550000 0.600000 ;
    END
  END sum_out[12]
  PIN sum_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 248.450000 0.000000 248.550000 0.600000 ;
    END
  END sum_out[11]
  PIN sum_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 247.450000 0.000000 247.550000 0.600000 ;
    END
  END sum_out[10]
  PIN sum_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 246.450000 0.000000 246.550000 0.600000 ;
    END
  END sum_out[9]
  PIN sum_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 245.450000 0.000000 245.550000 0.600000 ;
    END
  END sum_out[8]
  PIN sum_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 244.450000 0.000000 244.550000 0.600000 ;
    END
  END sum_out[7]
  PIN sum_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 243.450000 0.000000 243.550000 0.600000 ;
    END
  END sum_out[6]
  PIN sum_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 242.450000 0.000000 242.550000 0.600000 ;
    END
  END sum_out[5]
  PIN sum_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 241.450000 0.000000 241.550000 0.600000 ;
    END
  END sum_out[4]
  PIN sum_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 240.450000 0.000000 240.550000 0.600000 ;
    END
  END sum_out[3]
  PIN sum_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 239.450000 0.000000 239.550000 0.600000 ;
    END
  END sum_out[2]
  PIN sum_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 238.450000 0.000000 238.550000 0.600000 ;
    END
  END sum_out[1]
  PIN sum_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 237.450000 0.000000 237.550000 0.600000 ;
    END
  END sum_out[0]
  OBS
    LAYER M1 ;
      RECT 0.000000 0.000000 394.600000 394.400000 ;
    LAYER M2 ;
      RECT 0.000000 0.000000 394.600000 394.400000 ;
    LAYER M3 ;
      RECT 0.000000 243.150000 394.600000 394.400000 ;
      RECT 0.720000 242.850000 394.600000 243.150000 ;
      RECT 0.000000 242.150000 394.600000 242.850000 ;
      RECT 0.720000 241.850000 394.600000 242.150000 ;
      RECT 0.000000 241.150000 394.600000 241.850000 ;
      RECT 0.720000 240.850000 394.600000 241.150000 ;
      RECT 0.000000 240.150000 394.600000 240.850000 ;
      RECT 0.720000 239.850000 394.600000 240.150000 ;
      RECT 0.000000 239.150000 394.600000 239.850000 ;
      RECT 0.720000 238.850000 394.600000 239.150000 ;
      RECT 0.000000 238.150000 394.600000 238.850000 ;
      RECT 0.720000 237.850000 394.600000 238.150000 ;
      RECT 0.000000 237.150000 394.600000 237.850000 ;
      RECT 0.720000 236.850000 394.600000 237.150000 ;
      RECT 0.000000 236.150000 394.600000 236.850000 ;
      RECT 0.720000 235.850000 394.600000 236.150000 ;
      RECT 0.000000 235.150000 394.600000 235.850000 ;
      RECT 0.720000 234.850000 394.600000 235.150000 ;
      RECT 0.000000 234.150000 394.600000 234.850000 ;
      RECT 0.720000 233.850000 394.600000 234.150000 ;
      RECT 0.000000 233.150000 394.600000 233.850000 ;
      RECT 0.720000 232.850000 394.600000 233.150000 ;
      RECT 0.000000 232.150000 394.600000 232.850000 ;
      RECT 0.720000 231.850000 394.600000 232.150000 ;
      RECT 0.000000 231.150000 394.600000 231.850000 ;
      RECT 0.720000 230.850000 394.600000 231.150000 ;
      RECT 0.000000 230.150000 394.600000 230.850000 ;
      RECT 0.720000 229.850000 394.600000 230.150000 ;
      RECT 0.000000 229.150000 394.600000 229.850000 ;
      RECT 0.720000 228.850000 394.600000 229.150000 ;
      RECT 0.000000 228.150000 394.600000 228.850000 ;
      RECT 0.720000 227.850000 394.600000 228.150000 ;
      RECT 0.000000 227.150000 394.600000 227.850000 ;
      RECT 0.720000 226.850000 394.600000 227.150000 ;
      RECT 0.000000 226.150000 394.600000 226.850000 ;
      RECT 0.720000 225.850000 394.600000 226.150000 ;
      RECT 0.000000 225.150000 394.600000 225.850000 ;
      RECT 0.720000 224.850000 394.600000 225.150000 ;
      RECT 0.000000 224.150000 394.600000 224.850000 ;
      RECT 0.720000 223.850000 394.600000 224.150000 ;
      RECT 0.000000 223.150000 394.600000 223.850000 ;
      RECT 0.720000 222.850000 394.600000 223.150000 ;
      RECT 0.000000 222.150000 394.600000 222.850000 ;
      RECT 0.720000 221.850000 394.600000 222.150000 ;
      RECT 0.000000 221.150000 394.600000 221.850000 ;
      RECT 0.720000 220.850000 394.600000 221.150000 ;
      RECT 0.000000 220.150000 394.600000 220.850000 ;
      RECT 0.720000 219.850000 394.600000 220.150000 ;
      RECT 0.000000 219.150000 394.600000 219.850000 ;
      RECT 0.720000 218.850000 394.600000 219.150000 ;
      RECT 0.000000 218.150000 394.600000 218.850000 ;
      RECT 0.720000 217.850000 394.600000 218.150000 ;
      RECT 0.000000 217.150000 394.600000 217.850000 ;
      RECT 0.720000 216.850000 394.600000 217.150000 ;
      RECT 0.000000 216.150000 394.600000 216.850000 ;
      RECT 0.720000 215.850000 394.600000 216.150000 ;
      RECT 0.000000 215.150000 394.600000 215.850000 ;
      RECT 0.720000 214.850000 394.600000 215.150000 ;
      RECT 0.000000 214.150000 394.600000 214.850000 ;
      RECT 0.720000 213.850000 394.600000 214.150000 ;
      RECT 0.000000 213.150000 394.600000 213.850000 ;
      RECT 0.720000 212.850000 394.600000 213.150000 ;
      RECT 0.000000 212.150000 394.600000 212.850000 ;
      RECT 0.720000 211.850000 394.600000 212.150000 ;
      RECT 0.000000 211.150000 394.600000 211.850000 ;
      RECT 0.720000 210.850000 394.600000 211.150000 ;
      RECT 0.000000 210.150000 394.600000 210.850000 ;
      RECT 0.720000 209.850000 394.600000 210.150000 ;
      RECT 0.000000 209.150000 394.600000 209.850000 ;
      RECT 0.720000 208.850000 394.600000 209.150000 ;
      RECT 0.000000 208.150000 394.600000 208.850000 ;
      RECT 0.720000 207.850000 394.600000 208.150000 ;
      RECT 0.000000 207.150000 394.600000 207.850000 ;
      RECT 0.720000 206.850000 394.600000 207.150000 ;
      RECT 0.000000 206.150000 394.600000 206.850000 ;
      RECT 0.720000 205.850000 394.600000 206.150000 ;
      RECT 0.000000 205.150000 394.600000 205.850000 ;
      RECT 0.720000 204.850000 394.600000 205.150000 ;
      RECT 0.000000 204.150000 394.600000 204.850000 ;
      RECT 0.720000 203.850000 394.600000 204.150000 ;
      RECT 0.000000 203.150000 394.600000 203.850000 ;
      RECT 0.720000 202.850000 394.600000 203.150000 ;
      RECT 0.000000 202.150000 394.600000 202.850000 ;
      RECT 0.720000 201.850000 394.600000 202.150000 ;
      RECT 0.000000 201.150000 394.600000 201.850000 ;
      RECT 0.720000 200.850000 394.600000 201.150000 ;
      RECT 0.000000 200.150000 394.600000 200.850000 ;
      RECT 0.720000 199.850000 394.600000 200.150000 ;
      RECT 0.000000 199.150000 394.600000 199.850000 ;
      RECT 0.720000 198.850000 394.600000 199.150000 ;
      RECT 0.000000 198.150000 394.600000 198.850000 ;
      RECT 0.720000 197.850000 394.600000 198.150000 ;
      RECT 0.000000 197.150000 394.600000 197.850000 ;
      RECT 0.720000 196.850000 394.600000 197.150000 ;
      RECT 0.000000 196.150000 394.600000 196.850000 ;
      RECT 0.720000 195.850000 394.600000 196.150000 ;
      RECT 0.000000 195.150000 394.600000 195.850000 ;
      RECT 0.720000 194.850000 394.600000 195.150000 ;
      RECT 0.000000 194.150000 394.600000 194.850000 ;
      RECT 0.720000 193.850000 394.600000 194.150000 ;
      RECT 0.000000 193.150000 394.600000 193.850000 ;
      RECT 0.720000 192.850000 394.600000 193.150000 ;
      RECT 0.000000 192.150000 394.600000 192.850000 ;
      RECT 0.720000 191.850000 394.600000 192.150000 ;
      RECT 0.000000 191.150000 394.600000 191.850000 ;
      RECT 0.720000 190.850000 394.600000 191.150000 ;
      RECT 0.000000 190.150000 394.600000 190.850000 ;
      RECT 0.720000 189.850000 394.600000 190.150000 ;
      RECT 0.000000 189.150000 394.600000 189.850000 ;
      RECT 0.720000 188.850000 394.600000 189.150000 ;
      RECT 0.000000 188.150000 394.600000 188.850000 ;
      RECT 0.720000 187.850000 394.600000 188.150000 ;
      RECT 0.000000 187.150000 394.600000 187.850000 ;
      RECT 0.720000 186.850000 394.600000 187.150000 ;
      RECT 0.000000 186.150000 394.600000 186.850000 ;
      RECT 0.720000 185.850000 394.600000 186.150000 ;
      RECT 0.000000 185.150000 394.600000 185.850000 ;
      RECT 0.720000 184.850000 394.600000 185.150000 ;
      RECT 0.000000 184.150000 394.600000 184.850000 ;
      RECT 0.720000 183.850000 394.600000 184.150000 ;
      RECT 0.000000 183.150000 394.600000 183.850000 ;
      RECT 0.720000 182.850000 394.600000 183.150000 ;
      RECT 0.000000 182.150000 394.600000 182.850000 ;
      RECT 0.720000 181.850000 394.600000 182.150000 ;
      RECT 0.000000 181.150000 394.600000 181.850000 ;
      RECT 0.720000 180.850000 394.600000 181.150000 ;
      RECT 0.000000 180.150000 394.600000 180.850000 ;
      RECT 0.720000 179.850000 394.600000 180.150000 ;
      RECT 0.000000 179.150000 394.600000 179.850000 ;
      RECT 0.720000 178.850000 394.600000 179.150000 ;
      RECT 0.000000 178.150000 394.600000 178.850000 ;
      RECT 0.720000 177.850000 394.600000 178.150000 ;
      RECT 0.000000 177.150000 394.600000 177.850000 ;
      RECT 0.720000 176.850000 394.600000 177.150000 ;
      RECT 0.000000 176.150000 394.600000 176.850000 ;
      RECT 0.720000 175.850000 394.600000 176.150000 ;
      RECT 0.000000 175.150000 394.600000 175.850000 ;
      RECT 0.720000 174.850000 394.600000 175.150000 ;
      RECT 0.000000 174.150000 394.600000 174.850000 ;
      RECT 0.720000 173.850000 394.600000 174.150000 ;
      RECT 0.000000 173.150000 394.600000 173.850000 ;
      RECT 0.720000 172.850000 394.600000 173.150000 ;
      RECT 0.000000 172.150000 394.600000 172.850000 ;
      RECT 0.720000 171.850000 394.600000 172.150000 ;
      RECT 0.000000 171.150000 394.600000 171.850000 ;
      RECT 0.720000 170.850000 394.600000 171.150000 ;
      RECT 0.000000 170.150000 394.600000 170.850000 ;
      RECT 0.720000 169.850000 394.600000 170.150000 ;
      RECT 0.000000 169.150000 394.600000 169.850000 ;
      RECT 0.720000 168.850000 394.600000 169.150000 ;
      RECT 0.000000 168.150000 394.600000 168.850000 ;
      RECT 0.720000 167.850000 394.600000 168.150000 ;
      RECT 0.000000 167.150000 394.600000 167.850000 ;
      RECT 0.720000 166.850000 394.600000 167.150000 ;
      RECT 0.000000 166.150000 394.600000 166.850000 ;
      RECT 0.720000 165.850000 394.600000 166.150000 ;
      RECT 0.000000 165.150000 394.600000 165.850000 ;
      RECT 0.720000 164.850000 394.600000 165.150000 ;
      RECT 0.000000 164.150000 394.600000 164.850000 ;
      RECT 0.720000 163.850000 394.600000 164.150000 ;
      RECT 0.000000 163.150000 394.600000 163.850000 ;
      RECT 0.720000 162.850000 394.600000 163.150000 ;
      RECT 0.000000 162.150000 394.600000 162.850000 ;
      RECT 0.720000 161.850000 394.600000 162.150000 ;
      RECT 0.000000 161.150000 394.600000 161.850000 ;
      RECT 0.720000 160.850000 394.600000 161.150000 ;
      RECT 0.000000 160.150000 394.600000 160.850000 ;
      RECT 0.720000 159.850000 394.600000 160.150000 ;
      RECT 0.000000 159.150000 394.600000 159.850000 ;
      RECT 0.720000 158.850000 394.600000 159.150000 ;
      RECT 0.000000 158.150000 394.600000 158.850000 ;
      RECT 0.720000 157.850000 394.600000 158.150000 ;
      RECT 0.000000 157.150000 394.600000 157.850000 ;
      RECT 0.720000 156.850000 394.600000 157.150000 ;
      RECT 0.000000 156.150000 394.600000 156.850000 ;
      RECT 0.720000 155.850000 394.600000 156.150000 ;
      RECT 0.000000 155.150000 394.600000 155.850000 ;
      RECT 0.720000 154.850000 394.600000 155.150000 ;
      RECT 0.000000 154.150000 394.600000 154.850000 ;
      RECT 0.720000 153.850000 394.600000 154.150000 ;
      RECT 0.000000 153.150000 394.600000 153.850000 ;
      RECT 0.720000 152.850000 394.600000 153.150000 ;
      RECT 0.000000 152.150000 394.600000 152.850000 ;
      RECT 0.720000 151.850000 394.600000 152.150000 ;
      RECT 0.000000 151.150000 394.600000 151.850000 ;
      RECT 0.720000 150.850000 394.600000 151.150000 ;
      RECT 0.000000 0.760000 394.600000 150.850000 ;
      RECT 252.710000 0.000000 394.600000 0.760000 ;
      RECT 251.710000 0.000000 252.290000 0.760000 ;
      RECT 250.710000 0.000000 251.290000 0.760000 ;
      RECT 249.710000 0.000000 250.290000 0.760000 ;
      RECT 248.710000 0.000000 249.290000 0.760000 ;
      RECT 247.710000 0.000000 248.290000 0.760000 ;
      RECT 246.710000 0.000000 247.290000 0.760000 ;
      RECT 245.710000 0.000000 246.290000 0.760000 ;
      RECT 244.710000 0.000000 245.290000 0.760000 ;
      RECT 243.710000 0.000000 244.290000 0.760000 ;
      RECT 242.710000 0.000000 243.290000 0.760000 ;
      RECT 241.710000 0.000000 242.290000 0.760000 ;
      RECT 240.710000 0.000000 241.290000 0.760000 ;
      RECT 239.710000 0.000000 240.290000 0.760000 ;
      RECT 238.710000 0.000000 239.290000 0.760000 ;
      RECT 237.710000 0.000000 238.290000 0.760000 ;
      RECT 236.710000 0.000000 237.290000 0.760000 ;
      RECT 235.710000 0.000000 236.290000 0.760000 ;
      RECT 234.710000 0.000000 235.290000 0.760000 ;
      RECT 233.710000 0.000000 234.290000 0.760000 ;
      RECT 232.710000 0.000000 233.290000 0.760000 ;
      RECT 231.710000 0.000000 232.290000 0.760000 ;
      RECT 230.710000 0.000000 231.290000 0.760000 ;
      RECT 229.710000 0.000000 230.290000 0.760000 ;
      RECT 228.710000 0.000000 229.290000 0.760000 ;
      RECT 227.710000 0.000000 228.290000 0.760000 ;
      RECT 226.710000 0.000000 227.290000 0.760000 ;
      RECT 225.710000 0.000000 226.290000 0.760000 ;
      RECT 224.710000 0.000000 225.290000 0.760000 ;
      RECT 223.710000 0.000000 224.290000 0.760000 ;
      RECT 222.710000 0.000000 223.290000 0.760000 ;
      RECT 221.710000 0.000000 222.290000 0.760000 ;
      RECT 220.710000 0.000000 221.290000 0.760000 ;
      RECT 219.710000 0.000000 220.290000 0.760000 ;
      RECT 218.710000 0.000000 219.290000 0.760000 ;
      RECT 217.710000 0.000000 218.290000 0.760000 ;
      RECT 216.710000 0.000000 217.290000 0.760000 ;
      RECT 215.710000 0.000000 216.290000 0.760000 ;
      RECT 214.710000 0.000000 215.290000 0.760000 ;
      RECT 213.710000 0.000000 214.290000 0.760000 ;
      RECT 212.710000 0.000000 213.290000 0.760000 ;
      RECT 211.710000 0.000000 212.290000 0.760000 ;
      RECT 210.710000 0.000000 211.290000 0.760000 ;
      RECT 209.710000 0.000000 210.290000 0.760000 ;
      RECT 208.710000 0.000000 209.290000 0.760000 ;
      RECT 207.710000 0.000000 208.290000 0.760000 ;
      RECT 206.710000 0.000000 207.290000 0.760000 ;
      RECT 205.710000 0.000000 206.290000 0.760000 ;
      RECT 204.710000 0.000000 205.290000 0.760000 ;
      RECT 203.710000 0.000000 204.290000 0.760000 ;
      RECT 202.710000 0.000000 203.290000 0.760000 ;
      RECT 201.710000 0.000000 202.290000 0.760000 ;
      RECT 200.710000 0.000000 201.290000 0.760000 ;
      RECT 199.710000 0.000000 200.290000 0.760000 ;
      RECT 198.710000 0.000000 199.290000 0.760000 ;
      RECT 197.710000 0.000000 198.290000 0.760000 ;
      RECT 196.710000 0.000000 197.290000 0.760000 ;
      RECT 195.710000 0.000000 196.290000 0.760000 ;
      RECT 194.710000 0.000000 195.290000 0.760000 ;
      RECT 193.710000 0.000000 194.290000 0.760000 ;
      RECT 192.710000 0.000000 193.290000 0.760000 ;
      RECT 191.710000 0.000000 192.290000 0.760000 ;
      RECT 190.710000 0.000000 191.290000 0.760000 ;
      RECT 189.710000 0.000000 190.290000 0.760000 ;
      RECT 188.710000 0.000000 189.290000 0.760000 ;
      RECT 187.710000 0.000000 188.290000 0.760000 ;
      RECT 186.710000 0.000000 187.290000 0.760000 ;
      RECT 185.710000 0.000000 186.290000 0.760000 ;
      RECT 184.710000 0.000000 185.290000 0.760000 ;
      RECT 183.710000 0.000000 184.290000 0.760000 ;
      RECT 182.710000 0.000000 183.290000 0.760000 ;
      RECT 181.710000 0.000000 182.290000 0.760000 ;
      RECT 180.710000 0.000000 181.290000 0.760000 ;
      RECT 179.710000 0.000000 180.290000 0.760000 ;
      RECT 178.710000 0.000000 179.290000 0.760000 ;
      RECT 177.710000 0.000000 178.290000 0.760000 ;
      RECT 176.710000 0.000000 177.290000 0.760000 ;
      RECT 175.710000 0.000000 176.290000 0.760000 ;
      RECT 174.710000 0.000000 175.290000 0.760000 ;
      RECT 173.710000 0.000000 174.290000 0.760000 ;
      RECT 172.710000 0.000000 173.290000 0.760000 ;
      RECT 171.710000 0.000000 172.290000 0.760000 ;
      RECT 170.710000 0.000000 171.290000 0.760000 ;
      RECT 169.710000 0.000000 170.290000 0.760000 ;
      RECT 168.710000 0.000000 169.290000 0.760000 ;
      RECT 167.710000 0.000000 168.290000 0.760000 ;
      RECT 166.710000 0.000000 167.290000 0.760000 ;
      RECT 165.710000 0.000000 166.290000 0.760000 ;
      RECT 164.710000 0.000000 165.290000 0.760000 ;
      RECT 163.710000 0.000000 164.290000 0.760000 ;
      RECT 162.710000 0.000000 163.290000 0.760000 ;
      RECT 161.710000 0.000000 162.290000 0.760000 ;
      RECT 160.710000 0.000000 161.290000 0.760000 ;
      RECT 159.710000 0.000000 160.290000 0.760000 ;
      RECT 158.710000 0.000000 159.290000 0.760000 ;
      RECT 157.710000 0.000000 158.290000 0.760000 ;
      RECT 156.710000 0.000000 157.290000 0.760000 ;
      RECT 155.710000 0.000000 156.290000 0.760000 ;
      RECT 154.710000 0.000000 155.290000 0.760000 ;
      RECT 153.710000 0.000000 154.290000 0.760000 ;
      RECT 152.710000 0.000000 153.290000 0.760000 ;
      RECT 151.710000 0.000000 152.290000 0.760000 ;
      RECT 150.710000 0.000000 151.290000 0.760000 ;
      RECT 149.710000 0.000000 150.290000 0.760000 ;
      RECT 148.710000 0.000000 149.290000 0.760000 ;
      RECT 147.710000 0.000000 148.290000 0.760000 ;
      RECT 146.710000 0.000000 147.290000 0.760000 ;
      RECT 145.710000 0.000000 146.290000 0.760000 ;
      RECT 144.710000 0.000000 145.290000 0.760000 ;
      RECT 143.710000 0.000000 144.290000 0.760000 ;
      RECT 142.710000 0.000000 143.290000 0.760000 ;
      RECT 141.710000 0.000000 142.290000 0.760000 ;
      RECT 0.000000 0.000000 141.290000 0.760000 ;
    LAYER M4 ;
      RECT 0.000000 0.000000 394.600000 394.400000 ;
    LAYER M5 ;
      RECT 0.000000 0.000000 394.600000 394.400000 ;
    LAYER M6 ;
      RECT 0.000000 0.000000 394.600000 394.400000 ;
    LAYER M7 ;
      RECT 0.000000 0.000000 394.600000 394.400000 ;
    LAYER M8 ;
      RECT 0.000000 0.000000 394.600000 394.400000 ;
  END
END fullchip

END LIBRARY
